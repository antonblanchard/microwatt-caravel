
/* JTAG */
`include "tap_top.v"

/* UART */
`include "raminfr.v"
`include "uart_receiver.v"
`include "uart_rfifo.v"
`include "uart_tfifo.v"
`include "uart_transmitter.v"
`include "uart_defines.v"
`include "uart_regs.v"
`include "uart_sync_flops.v"
`include "uart_wb.v"
`include "uart_top.v"
`include "simplebus_host.v"
module plru_1
  (input  clk,
   input  rst,
   input  acc,
   input  acc_en,
   output lru);
  wire [1:0] tree;
  wire n33606_o;
  wire n33613_o;
  wire n33614_o;
  wire n33615_o;
  wire n33620_o;
  wire n33621_o;
  wire n33623_o;
  wire [1:0] n33626_o;
  reg [1:0] n33633_q;
  assign lru = n33606_o;
  /* plru.vhdl:26:12  */
  assign tree = n33633_q; // (signal)
  /* plru.vhdl:38:34  */
  assign n33606_o = tree[1];
  /* plru.vhdl:61:35  */
  assign n33613_o = ~acc;
  assign n33614_o = tree[1];
  /* plru.vhdl:57:13  */
  assign n33615_o = acc_en ? n33613_o : n33614_o;
  assign n33620_o = tree[0];
  /* plru.vhdl:55:13  */
  assign n33621_o = rst ? 1'b0 : n33620_o;
  /* plru.vhdl:55:13  */
  assign n33623_o = rst ? 1'b0 : n33615_o;
  assign n33626_o = {n33623_o, n33621_o};
  /* plru.vhdl:54:9  */
  always @(posedge clk)
    n33633_q <= n33626_o;
endmodule

module pmu
  (input  clk,
   input  rst,
   input  p_in_mfspr,
   input  p_in_mtspr,
   input  [4:0] p_in_spr_num,
   input  [63:0] p_in_spr_val,
   input  [3:0] p_in_tbbits,
   input  p_in_pmm_msr,
   input  p_in_pr_msr,
   input  p_in_run,
   input  [63:0] p_in_nia,
   input  [63:0] p_in_addr,
   input  p_in_addr_v,
   input  [20:0] p_in_occur,
   output [63:0] p_out_spr_val,
   output p_out_intr);
  wire [227:0] n32886_o;
  wire [63:0] n32888_o;
  wire n32889_o;
  wire [191:0] pmcs;
  wire [31:0] mmcr0;
  wire [63:0] mmcr1;
  wire [63:0] mmcr2;
  wire [63:0] mmcra;
  wire [63:0] siar;
  wire [63:0] sdar;
  wire [63:0] sier;
  wire [5:0] doinc;
  wire doalert;
  wire doevent;
  wire [3:0] prev_tb;
  wire [3:0] n32890_o;
  wire [31:0] n32891_o;
  wire [63:0] n32893_o;
  wire n32895_o;
  wire [31:0] n32896_o;
  wire [63:0] n32898_o;
  wire n32900_o;
  wire [31:0] n32901_o;
  wire [63:0] n32903_o;
  wire n32905_o;
  wire [31:0] n32906_o;
  wire [63:0] n32908_o;
  wire n32910_o;
  wire [31:0] n32911_o;
  wire [63:0] n32913_o;
  wire n32915_o;
  wire [31:0] n32916_o;
  wire [63:0] n32918_o;
  wire n32920_o;
  wire [63:0] n32922_o;
  wire n32924_o;
  wire n32926_o;
  wire n32928_o;
  wire n32930_o;
  wire n32932_o;
  wire n32934_o;
  wire n32936_o;
  wire [12:0] n32938_o;
  reg [63:0] n32939_o;
  wire n32940_o;
  wire n32943_o;
  wire [3:0] n32944_o;
  wire [30:0] n32945_o;
  wire [31:0] n32946_o;
  wire n32948_o;
  wire n32949_o;
  wire [31:0] n32950_o;
  wire n32951_o;
  wire [31:0] n32952_o;
  wire [31:0] n32954_o;
  wire [31:0] n32955_o;
  wire [31:0] n32956_o;
  wire [31:0] n32957_o;
  wire n32958_o;
  wire [3:0] n32959_o;
  wire [30:0] n32960_o;
  wire [31:0] n32961_o;
  wire n32963_o;
  wire n32964_o;
  wire [31:0] n32965_o;
  wire n32966_o;
  wire [31:0] n32967_o;
  wire [31:0] n32969_o;
  wire [31:0] n32970_o;
  wire [31:0] n32971_o;
  wire [31:0] n32972_o;
  wire n32973_o;
  wire [3:0] n32974_o;
  wire [30:0] n32975_o;
  wire [31:0] n32976_o;
  wire n32978_o;
  wire n32979_o;
  wire [31:0] n32980_o;
  wire n32981_o;
  wire [31:0] n32982_o;
  wire [31:0] n32984_o;
  wire [31:0] n32985_o;
  wire [31:0] n32986_o;
  wire [31:0] n32987_o;
  wire n32988_o;
  wire [3:0] n32989_o;
  wire [30:0] n32990_o;
  wire [31:0] n32991_o;
  wire n32993_o;
  wire n32994_o;
  wire [31:0] n32995_o;
  wire n32996_o;
  wire [31:0] n32997_o;
  wire [31:0] n32999_o;
  wire [31:0] n33000_o;
  wire [31:0] n33001_o;
  wire [31:0] n33002_o;
  wire n33003_o;
  wire [3:0] n33004_o;
  wire [30:0] n33005_o;
  wire [31:0] n33006_o;
  wire n33008_o;
  wire n33009_o;
  wire [31:0] n33010_o;
  wire n33011_o;
  wire [31:0] n33012_o;
  wire [31:0] n33014_o;
  wire [31:0] n33015_o;
  wire [31:0] n33016_o;
  wire [31:0] n33017_o;
  wire n33018_o;
  wire [3:0] n33019_o;
  wire [30:0] n33020_o;
  wire [31:0] n33021_o;
  wire n33023_o;
  wire n33024_o;
  wire [31:0] n33025_o;
  wire n33026_o;
  wire [31:0] n33027_o;
  wire [31:0] n33029_o;
  wire [31:0] n33030_o;
  wire [31:0] n33031_o;
  wire [31:0] n33032_o;
  wire n33033_o;
  wire [3:0] n33034_o;
  wire n33036_o;
  wire n33037_o;
  wire [9:0] n33040_o;
  wire [19:0] n33043_o;
  wire n33047_o;
  wire n33048_o;
  wire n33049_o;
  wire n33050_o;
  wire n33051_o;
  wire n33052_o;
  wire n33053_o;
  wire n33054_o;
  wire n33055_o;
  wire n33056_o;
  wire n33057_o;
  wire n33059_o;
  wire n33060_o;
  wire n33061_o;
  wire n33062_o;
  wire n33063_o;
  wire n33064_o;
  wire n33066_o;
  wire n33067_o;
  wire [31:0] n33068_o;
  wire [6:0] n33069_o;
  wire [6:0] n33070_o;
  wire [6:0] n33071_o;
  wire n33072_o;
  wire n33073_o;
  wire [2:0] n33074_o;
  wire [2:0] n33075_o;
  wire [2:0] n33076_o;
  wire n33077_o;
  wire n33078_o;
  wire n33079_o;
  wire n33080_o;
  wire n33081_o;
  wire n33082_o;
  wire n33083_o;
  wire [11:0] n33084_o;
  wire [11:0] n33085_o;
  wire [11:0] n33086_o;
  wire n33087_o;
  wire n33088_o;
  wire [3:0] n33089_o;
  wire [3:0] n33090_o;
  wire [3:0] n33091_o;
  wire n33092_o;
  wire n33093_o;
  wire n33094_o;
  wire [3:0] n33095_o;
  wire n33097_o;
  wire n33098_o;
  wire [63:0] n33099_o;
  wire [63:0] n33100_o;
  wire n33101_o;
  wire [3:0] n33102_o;
  wire n33104_o;
  wire n33105_o;
  wire [63:0] n33106_o;
  wire [63:0] n33107_o;
  wire n33108_o;
  wire [3:0] n33109_o;
  wire n33111_o;
  wire n33112_o;
  wire [62:0] n33115_o;
  wire [63:0] n33116_o;
  wire [63:0] n33117_o;
  wire n33118_o;
  wire [3:0] n33119_o;
  wire n33121_o;
  wire n33122_o;
  wire [63:0] n33123_o;
  wire [63:0] n33124_o;
  wire [63:0] n33125_o;
  wire [63:0] n33126_o;
  wire n33127_o;
  wire [3:0] n33128_o;
  wire n33130_o;
  wire n33131_o;
  wire [63:0] n33132_o;
  wire [63:0] n33133_o;
  wire [63:0] n33134_o;
  wire [63:0] n33135_o;
  wire n33136_o;
  wire [3:0] n33137_o;
  wire n33139_o;
  wire n33140_o;
  wire [63:0] n33141_o;
  wire n33142_o;
  localparam [63:0] n33143_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire [37:0] n33144_o;
  wire [1:0] n33147_o;
  wire n33149_o;
  wire [20:0] n33150_o;
  wire [63:0] n33151_o;
  wire [63:0] n33152_o;
  wire [63:0] n33153_o;
  wire [191:0] n33154_o;
  wire [191:0] n33155_o;
  wire [31:0] n33156_o;
  wire [31:0] n33158_o;
  wire [63:0] n33159_o;
  wire [63:0] n33160_o;
  wire [63:0] n33161_o;
  wire [63:0] n33162_o;
  wire [63:0] n33163_o;
  wire [63:0] n33164_o;
  wire [3:0] n33165_o;
  wire [3:0] n33184_o;
  wire [3:0] n33185_o;
  wire [3:0] n33186_o;
  wire [1:0] n33187_o;
  wire [30:0] n33188_o;
  wire [31:0] n33189_o;
  wire [31:0] n33191_o;
  wire [1:0] n33192_o;
  wire n33195_o;
  wire n33196_o;
  wire n33199_o;
  wire n33201_o;
  wire n33202_o;
  wire n33203_o;
  wire n33205_o;
  wire n33206_o;
  wire n33207_o;
  wire n33208_o;
  wire n33209_o;
  wire n33210_o;
  wire n33211_o;
  wire n33212_o;
  wire n33214_o;
  wire n33215_o;
  wire [1:0] n33216_o;
  wire n33218_o;
  wire n33219_o;
  wire n33220_o;
  wire n33221_o;
  wire n33222_o;
  wire n33223_o;
  wire n33225_o;
  wire [7:0] n33226_o;
  wire n33229_o;
  wire [20:0] n33230_o;
  wire n33231_o;
  wire n33233_o;
  wire n33235_o;
  wire n33236_o;
  wire [20:0] n33237_o;
  wire n33238_o;
  wire n33240_o;
  wire [20:0] n33241_o;
  wire n33242_o;
  wire n33244_o;
  wire [20:0] n33245_o;
  wire n33246_o;
  wire n33248_o;
  wire n33249_o;
  wire n33251_o;
  wire [20:0] n33252_o;
  wire n33253_o;
  wire n33255_o;
  wire [6:0] n33256_o;
  reg n33258_o;
  localparam [5:0] n33259_o = 6'b000000;
  reg n33263_o;
  wire [7:0] n33265_o;
  wire [20:0] n33266_o;
  wire n33267_o;
  wire n33269_o;
  wire [20:0] n33270_o;
  wire n33271_o;
  wire n33273_o;
  wire n33274_o;
  wire n33276_o;
  wire [20:0] n33277_o;
  wire n33278_o;
  wire n33280_o;
  wire [20:0] n33281_o;
  wire n33282_o;
  wire n33284_o;
  wire [20:0] n33285_o;
  wire n33286_o;
  wire n33288_o;
  wire [20:0] n33289_o;
  wire n33290_o;
  wire n33292_o;
  wire [20:0] n33293_o;
  wire n33294_o;
  wire n33296_o;
  wire [7:0] n33297_o;
  wire n33298_o;
  reg n33299_o;
  wire [7:0] n33301_o;
  wire [20:0] n33302_o;
  wire n33303_o;
  wire n33305_o;
  wire [20:0] n33306_o;
  wire n33307_o;
  wire n33309_o;
  wire [20:0] n33310_o;
  wire n33311_o;
  wire n33312_o;
  wire n33313_o;
  wire n33315_o;
  wire [20:0] n33316_o;
  wire n33317_o;
  wire n33319_o;
  wire n33321_o;
  wire [20:0] n33322_o;
  wire n33323_o;
  wire n33325_o;
  wire [5:0] n33326_o;
  wire n33327_o;
  reg n33328_o;
  wire [7:0] n33330_o;
  wire [20:0] n33331_o;
  wire n33332_o;
  wire n33334_o;
  wire [20:0] n33335_o;
  wire n33336_o;
  wire n33338_o;
  wire n33339_o;
  wire n33341_o;
  wire [20:0] n33342_o;
  wire n33343_o;
  wire n33345_o;
  wire [20:0] n33346_o;
  wire n33347_o;
  wire n33349_o;
  wire [20:0] n33350_o;
  wire n33351_o;
  wire n33352_o;
  wire n33353_o;
  wire n33355_o;
  wire [20:0] n33356_o;
  wire n33357_o;
  wire n33359_o;
  wire [20:0] n33360_o;
  wire n33361_o;
  wire n33363_o;
  wire [7:0] n33364_o;
  wire n33365_o;
  reg n33366_o;
  wire n33368_o;
  wire n33369_o;
  wire n33370_o;
  wire [20:0] n33371_o;
  wire n33372_o;
  wire n33373_o;
  wire n33375_o;
  wire n33376_o;
  wire n33377_o;
  wire n33378_o;
  wire n33379_o;
  wire n33380_o;
  wire n33381_o;
  wire n33382_o;
  wire n33383_o;
  wire n33384_o;
  wire n33385_o;
  wire n33386_o;
  wire n33387_o;
  wire n33388_o;
  wire n33389_o;
  wire n33390_o;
  wire n33391_o;
  wire n33392_o;
  wire n33393_o;
  wire n33394_o;
  wire n33395_o;
  wire n33396_o;
  wire n33397_o;
  wire n33398_o;
  wire n33399_o;
  wire n33400_o;
  wire n33401_o;
  wire n33402_o;
  wire n33403_o;
  wire n33404_o;
  wire n33405_o;
  wire n33406_o;
  wire n33407_o;
  wire n33408_o;
  wire n33409_o;
  wire n33410_o;
  wire n33411_o;
  wire n33412_o;
  wire n33413_o;
  wire n33414_o;
  wire n33415_o;
  wire n33417_o;
  wire n33418_o;
  wire n33419_o;
  wire n33420_o;
  wire n33421_o;
  wire n33422_o;
  wire n33423_o;
  wire n33424_o;
  wire [2:0] n33426_o;
  wire [2:0] n33427_o;
  wire n33428_o;
  wire n33429_o;
  wire [1:0] n33431_o;
  wire [1:0] n33432_o;
  wire n33433_o;
  localparam [4:0] n33434_o = 5'b00000;
  wire [4:0] n33435_o;
  wire n33437_o;
  wire n33438_o;
  wire n33439_o;
  wire n33440_o;
  wire n33441_o;
  wire n33442_o;
  wire n33443_o;
  wire n33444_o;
  wire n33445_o;
  wire n33446_o;
  wire n33447_o;
  wire n33448_o;
  wire n33449_o;
  wire n33450_o;
  wire n33451_o;
  wire n33452_o;
  wire n33454_o;
  wire n33455_o;
  wire n33456_o;
  wire n33457_o;
  wire n33458_o;
  wire n33459_o;
  wire n33460_o;
  wire n33461_o;
  wire n33462_o;
  wire n33463_o;
  wire n33464_o;
  wire n33465_o;
  wire n33466_o;
  wire n33467_o;
  wire n33468_o;
  wire n33469_o;
  wire n33470_o;
  wire n33472_o;
  wire n33473_o;
  wire n33474_o;
  wire n33475_o;
  wire n33479_o;
  wire n33480_o;
  wire n33481_o;
  wire n33482_o;
  wire n33483_o;
  wire n33484_o;
  wire n33485_o;
  wire n33486_o;
  wire n33487_o;
  wire n33488_o;
  wire n33489_o;
  wire n33490_o;
  wire n33491_o;
  wire n33492_o;
  wire n33493_o;
  wire n33494_o;
  wire n33496_o;
  wire n33497_o;
  wire n33498_o;
  wire n33499_o;
  wire n33503_o;
  wire n33504_o;
  wire n33505_o;
  wire n33506_o;
  wire n33507_o;
  wire n33508_o;
  wire n33509_o;
  wire n33510_o;
  wire n33511_o;
  wire n33512_o;
  wire n33513_o;
  wire n33514_o;
  wire n33515_o;
  wire n33516_o;
  wire n33517_o;
  wire n33518_o;
  wire n33520_o;
  wire n33521_o;
  wire n33522_o;
  wire n33523_o;
  wire n33527_o;
  wire n33528_o;
  wire n33529_o;
  wire n33530_o;
  wire n33531_o;
  wire n33532_o;
  wire n33533_o;
  wire n33534_o;
  wire n33535_o;
  wire n33536_o;
  wire n33537_o;
  wire n33538_o;
  wire n33539_o;
  wire n33540_o;
  wire n33541_o;
  wire n33542_o;
  wire n33544_o;
  wire n33545_o;
  wire n33546_o;
  wire n33547_o;
  wire n33548_o;
  wire n33549_o;
  wire n33550_o;
  wire n33551_o;
  wire n33552_o;
  wire n33553_o;
  wire n33554_o;
  wire n33555_o;
  wire n33556_o;
  wire n33557_o;
  wire n33558_o;
  wire n33559_o;
  wire n33560_o;
  wire n33561_o;
  wire n33562_o;
  wire n33563_o;
  wire n33564_o;
  wire n33565_o;
  wire n33566_o;
  wire n33568_o;
  wire [1:0] n33569_o;
  wire n33571_o;
  wire n33572_o;
  wire [20:0] n33573_o;
  wire n33574_o;
  wire n33575_o;
  wire n33576_o;
  wire [1:0] n33577_o;
  wire [1:0] n33578_o;
  wire [1:0] n33579_o;
  wire [5:0] n33580_o;
  wire n33581_o;
  wire n33582_o;
  reg [191:0] n33587_q;
  reg [31:0] n33588_q;
  reg [63:0] n33589_q;
  reg [63:0] n33590_q;
  reg [63:0] n33591_q;
  reg [63:0] n33592_q;
  reg [63:0] n33593_q;
  reg [63:0] n33594_q;
  reg [3:0] n33595_q;
  wire [64:0] n33596_o;
  wire n33597_o;
  wire n33598_o;
  wire n33599_o;
  wire n33600_o;
  wire [1:0] n33601_o;
  reg n33602_o;
  assign p_out_spr_val = n32888_o;
  assign p_out_intr = n32889_o;
  /* nonrandom.vhdl:11:9  */
  assign n32886_o = {p_in_occur, p_in_addr_v, p_in_addr, p_in_nia, p_in_run, p_in_pr_msr, p_in_pmm_msr, p_in_tbbits, p_in_spr_val, p_in_spr_num, p_in_mtspr, p_in_mfspr};
  assign n32888_o = n33596_o[63:0];
  /* divider.vhdl:39:13  */
  assign n32889_o = n33596_o[64];
  /* pmu.vhdl:108:12  */
  assign pmcs = n33587_q; // (signal)
  /* pmu.vhdl:109:12  */
  assign mmcr0 = n33588_q; // (signal)
  /* pmu.vhdl:110:12  */
  assign mmcr1 = n33589_q; // (signal)
  /* pmu.vhdl:111:12  */
  assign mmcr2 = n33590_q; // (signal)
  /* pmu.vhdl:112:12  */
  assign mmcra = n33591_q; // (signal)
  /* pmu.vhdl:113:12  */
  assign siar = n33592_q; // (signal)
  /* pmu.vhdl:114:12  */
  assign sdar = n33593_q; // (signal)
  /* pmu.vhdl:115:12  */
  assign sier = n33594_q; // (signal)
  /* pmu.vhdl:117:12  */
  assign doinc = n33580_o; // (signal)
  /* pmu.vhdl:118:12  */
  assign doalert = n33582_o; // (signal)
  /* pmu.vhdl:119:12  */
  assign doevent = n33225_o; // (signal)
  /* pmu.vhdl:121:12  */
  assign prev_tb = n33595_q; // (signal)
  /* pmu.vhdl:125:22  */
  assign n32890_o = n32886_o[5:2];
  /* pmu.vhdl:126:22  */
  assign n32891_o = pmcs[191:160];
  /* pmu.vhdl:126:16  */
  assign n32893_o = {32'b00000000000000000000000000000000, n32891_o};
  /* pmu.vhdl:126:26  */
  assign n32895_o = n32890_o == 4'b0011;
  /* pmu.vhdl:127:22  */
  assign n32896_o = pmcs[159:128];
  /* pmu.vhdl:127:16  */
  assign n32898_o = {32'b00000000000000000000000000000000, n32896_o};
  /* pmu.vhdl:127:26  */
  assign n32900_o = n32890_o == 4'b0100;
  /* pmu.vhdl:128:22  */
  assign n32901_o = pmcs[127:96];
  /* pmu.vhdl:128:16  */
  assign n32903_o = {32'b00000000000000000000000000000000, n32901_o};
  /* pmu.vhdl:128:26  */
  assign n32905_o = n32890_o == 4'b0101;
  /* pmu.vhdl:129:22  */
  assign n32906_o = pmcs[95:64];
  /* pmu.vhdl:129:16  */
  assign n32908_o = {32'b00000000000000000000000000000000, n32906_o};
  /* pmu.vhdl:129:26  */
  assign n32910_o = n32890_o == 4'b0110;
  /* pmu.vhdl:130:22  */
  assign n32911_o = pmcs[63:32];
  /* pmu.vhdl:130:16  */
  assign n32913_o = {32'b00000000000000000000000000000000, n32911_o};
  /* pmu.vhdl:130:26  */
  assign n32915_o = n32890_o == 4'b0111;
  /* pmu.vhdl:131:22  */
  assign n32916_o = pmcs[31:0];
  /* pmu.vhdl:131:16  */
  assign n32918_o = {32'b00000000000000000000000000000000, n32916_o};
  /* pmu.vhdl:131:26  */
  assign n32920_o = n32890_o == 4'b1000;
  /* pmu.vhdl:132:16  */
  assign n32922_o = {32'b00000000000000000000000000000000, mmcr0};
  /* pmu.vhdl:132:26  */
  assign n32924_o = n32890_o == 4'b1011;
  /* pmu.vhdl:133:26  */
  assign n32926_o = n32890_o == 4'b1110;
  /* pmu.vhdl:134:26  */
  assign n32928_o = n32890_o == 4'b0001;
  /* pmu.vhdl:135:26  */
  assign n32930_o = n32890_o == 4'b0010;
  /* pmu.vhdl:136:26  */
  assign n32932_o = n32890_o == 4'b1100;
  /* pmu.vhdl:137:26  */
  assign n32934_o = n32890_o == 4'b1101;
  /* pmu.vhdl:138:26  */
  assign n32936_o = n32890_o == 4'b0000;
  assign n32938_o = {n32936_o, n32934_o, n32932_o, n32930_o, n32928_o, n32926_o, n32924_o, n32920_o, n32915_o, n32910_o, n32905_o, n32900_o, n32895_o};
  /* pmu.vhdl:125:5  */
  always @*
    case (n32938_o)
      13'b1000000000000: n32939_o = sier;
      13'b0100000000000: n32939_o = sdar;
      13'b0010000000000: n32939_o = siar;
      13'b0001000000000: n32939_o = mmcra;
      13'b0000100000000: n32939_o = mmcr2;
      13'b0000010000000: n32939_o = mmcr1;
      13'b0000001000000: n32939_o = n32922_o;
      13'b0000000100000: n32939_o = n32918_o;
      13'b0000000010000: n32939_o = n32913_o;
      13'b0000000001000: n32939_o = n32908_o;
      13'b0000000000100: n32939_o = n32903_o;
      13'b0000000000010: n32939_o = n32898_o;
      13'b0000000000001: n32939_o = n32893_o;
      default: n32939_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* pmu.vhdl:141:24  */
  assign n32940_o = mmcr0[7];
  /* pmu.vhdl:150:29  */
  assign n32943_o = n32886_o[1];
  /* pmu.vhdl:150:77  */
  assign n32944_o = n32886_o[5:2];
  /* pmu.vhdl:150:45  */
  assign n32945_o = {27'b0, n32944_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n32946_o = {1'b0, n32945_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n32948_o = n32946_o == 32'b00000000000000000000000000000011;
  /* pmu.vhdl:150:41  */
  assign n32949_o = n32943_o & n32948_o;
  /* pmu.vhdl:151:48  */
  assign n32950_o = n32886_o[38:7];
  /* pmu.vhdl:152:32  */
  assign n32951_o = doinc[5];
  /* pmu.vhdl:153:67  */
  assign n32952_o = pmcs[191:160];
  /* pmu.vhdl:153:72  */
  assign n32954_o = n32952_o + 32'b00000000000000000000000000000001;
  assign n32955_o = pmcs[191:160];
  /* pmu.vhdl:152:21  */
  assign n32956_o = n32951_o ? n32954_o : n32955_o;
  /* pmu.vhdl:150:21  */
  assign n32957_o = n32949_o ? n32950_o : n32956_o;
  /* pmu.vhdl:150:29  */
  assign n32958_o = n32886_o[1];
  /* pmu.vhdl:150:77  */
  assign n32959_o = n32886_o[5:2];
  /* pmu.vhdl:150:45  */
  assign n32960_o = {27'b0, n32959_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n32961_o = {1'b0, n32960_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n32963_o = n32961_o == 32'b00000000000000000000000000000100;
  /* pmu.vhdl:150:41  */
  assign n32964_o = n32958_o & n32963_o;
  /* pmu.vhdl:151:48  */
  assign n32965_o = n32886_o[38:7];
  /* pmu.vhdl:152:32  */
  assign n32966_o = doinc[4];
  /* pmu.vhdl:153:67  */
  assign n32967_o = pmcs[159:128];
  /* pmu.vhdl:153:72  */
  assign n32969_o = n32967_o + 32'b00000000000000000000000000000001;
  assign n32970_o = pmcs[159:128];
  /* pmu.vhdl:152:21  */
  assign n32971_o = n32966_o ? n32969_o : n32970_o;
  /* pmu.vhdl:150:21  */
  assign n32972_o = n32964_o ? n32965_o : n32971_o;
  /* pmu.vhdl:150:29  */
  assign n32973_o = n32886_o[1];
  /* pmu.vhdl:150:77  */
  assign n32974_o = n32886_o[5:2];
  /* pmu.vhdl:150:45  */
  assign n32975_o = {27'b0, n32974_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n32976_o = {1'b0, n32975_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n32978_o = n32976_o == 32'b00000000000000000000000000000101;
  /* pmu.vhdl:150:41  */
  assign n32979_o = n32973_o & n32978_o;
  /* pmu.vhdl:151:48  */
  assign n32980_o = n32886_o[38:7];
  /* pmu.vhdl:152:32  */
  assign n32981_o = doinc[3];
  /* pmu.vhdl:153:67  */
  assign n32982_o = pmcs[127:96];
  /* pmu.vhdl:153:72  */
  assign n32984_o = n32982_o + 32'b00000000000000000000000000000001;
  assign n32985_o = pmcs[127:96];
  /* pmu.vhdl:152:21  */
  assign n32986_o = n32981_o ? n32984_o : n32985_o;
  /* pmu.vhdl:150:21  */
  assign n32987_o = n32979_o ? n32980_o : n32986_o;
  /* pmu.vhdl:150:29  */
  assign n32988_o = n32886_o[1];
  /* pmu.vhdl:150:77  */
  assign n32989_o = n32886_o[5:2];
  /* pmu.vhdl:150:45  */
  assign n32990_o = {27'b0, n32989_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n32991_o = {1'b0, n32990_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n32993_o = n32991_o == 32'b00000000000000000000000000000110;
  /* pmu.vhdl:150:41  */
  assign n32994_o = n32988_o & n32993_o;
  /* pmu.vhdl:151:48  */
  assign n32995_o = n32886_o[38:7];
  /* pmu.vhdl:152:32  */
  assign n32996_o = doinc[2];
  /* pmu.vhdl:153:67  */
  assign n32997_o = pmcs[95:64];
  /* pmu.vhdl:153:72  */
  assign n32999_o = n32997_o + 32'b00000000000000000000000000000001;
  assign n33000_o = pmcs[95:64];
  /* pmu.vhdl:152:21  */
  assign n33001_o = n32996_o ? n32999_o : n33000_o;
  /* pmu.vhdl:150:21  */
  assign n33002_o = n32994_o ? n32995_o : n33001_o;
  /* pmu.vhdl:150:29  */
  assign n33003_o = n32886_o[1];
  /* pmu.vhdl:150:77  */
  assign n33004_o = n32886_o[5:2];
  /* pmu.vhdl:150:45  */
  assign n33005_o = {27'b0, n33004_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n33006_o = {1'b0, n33005_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n33008_o = n33006_o == 32'b00000000000000000000000000000111;
  /* pmu.vhdl:150:41  */
  assign n33009_o = n33003_o & n33008_o;
  /* pmu.vhdl:151:48  */
  assign n33010_o = n32886_o[38:7];
  /* pmu.vhdl:152:32  */
  assign n33011_o = doinc[1];
  /* pmu.vhdl:153:67  */
  assign n33012_o = pmcs[63:32];
  /* pmu.vhdl:153:72  */
  assign n33014_o = n33012_o + 32'b00000000000000000000000000000001;
  assign n33015_o = pmcs[63:32];
  /* pmu.vhdl:152:21  */
  assign n33016_o = n33011_o ? n33014_o : n33015_o;
  /* pmu.vhdl:150:21  */
  assign n33017_o = n33009_o ? n33010_o : n33016_o;
  /* pmu.vhdl:150:29  */
  assign n33018_o = n32886_o[1];
  /* pmu.vhdl:150:77  */
  assign n33019_o = n32886_o[5:2];
  /* pmu.vhdl:150:45  */
  assign n33020_o = {27'b0, n33019_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n33021_o = {1'b0, n33020_o};  //  uext
  /* pmu.vhdl:150:92  */
  assign n33023_o = n33021_o == 32'b00000000000000000000000000001000;
  /* pmu.vhdl:150:41  */
  assign n33024_o = n33018_o & n33023_o;
  /* pmu.vhdl:151:48  */
  assign n33025_o = n32886_o[38:7];
  /* pmu.vhdl:152:32  */
  assign n33026_o = doinc[0];
  /* pmu.vhdl:153:67  */
  assign n33027_o = pmcs[31:0];
  /* pmu.vhdl:153:72  */
  assign n33029_o = n33027_o + 32'b00000000000000000000000000000001;
  assign n33030_o = pmcs[31:0];
  /* pmu.vhdl:152:21  */
  assign n33031_o = n33026_o ? n33029_o : n33030_o;
  /* pmu.vhdl:150:21  */
  assign n33032_o = n33024_o ? n33025_o : n33031_o;
  /* pmu.vhdl:156:25  */
  assign n33033_o = n32886_o[1];
  /* pmu.vhdl:156:53  */
  assign n33034_o = n32886_o[5:2];
  /* pmu.vhdl:156:66  */
  assign n33036_o = n33034_o == 4'b1011;
  /* pmu.vhdl:156:37  */
  assign n33037_o = n33033_o & n33036_o;
  assign n33040_o = n32886_o[38:29];
  assign n33043_o = n32886_o[26:7];
  assign n33047_o = mmcr0[7];
  /* pmu.vhdl:161:21  */
  assign n33048_o = doalert ? 1'b1 : n33047_o;
  assign n33049_o = mmcr0[11];
  /* pmu.vhdl:161:21  */
  assign n33050_o = doalert ? 1'b0 : n33049_o;
  assign n33051_o = mmcr0[26];
  /* pmu.vhdl:161:21  */
  assign n33052_o = doalert ? 1'b0 : n33051_o;
  /* pmu.vhdl:166:47  */
  assign n33053_o = mmcr0[25];
  /* pmu.vhdl:166:38  */
  assign n33054_o = doevent & n33053_o;
  /* pmu.vhdl:166:76  */
  assign n33055_o = mmcr0[13];
  /* pmu.vhdl:166:92  */
  assign n33056_o = ~n33055_o;
  /* pmu.vhdl:166:67  */
  assign n33057_o = n33054_o & n33056_o;
  assign n33059_o = mmcr0[31];
  /* pmu.vhdl:166:21  */
  assign n33060_o = n33057_o ? 1'b1 : n33059_o;
  /* pmu.vhdl:169:49  */
  assign n33061_o = pmcs[191];
  /* pmu.vhdl:169:39  */
  assign n33062_o = doevent | n33061_o;
  /* pmu.vhdl:169:70  */
  assign n33063_o = mmcr0[13];
  /* pmu.vhdl:169:61  */
  assign n33064_o = n33062_o & n33063_o;
  assign n33066_o = mmcr0[13];
  /* pmu.vhdl:169:21  */
  assign n33067_o = n33064_o ? 1'b0 : n33066_o;
  assign n33068_o = {n33040_o, 1'b0, 1'b0, n33043_o};
  assign n33069_o = n33068_o[6:0];
  assign n33070_o = mmcr0[6:0];
  /* pmu.vhdl:156:17  */
  assign n33071_o = n33037_o ? n33069_o : n33070_o;
  assign n33072_o = n33068_o[7];
  /* pmu.vhdl:156:17  */
  assign n33073_o = n33037_o ? n33072_o : n33048_o;
  assign n33074_o = n33068_o[10:8];
  assign n33075_o = mmcr0[10:8];
  /* pmu.vhdl:156:17  */
  assign n33076_o = n33037_o ? n33074_o : n33075_o;
  assign n33077_o = n33068_o[11];
  /* pmu.vhdl:156:17  */
  assign n33078_o = n33037_o ? n33077_o : n33050_o;
  assign n33079_o = n33068_o[12];
  assign n33080_o = mmcr0[12];
  /* pmu.vhdl:156:17  */
  assign n33081_o = n33037_o ? n33079_o : n33080_o;
  assign n33082_o = n33068_o[13];
  /* pmu.vhdl:156:17  */
  assign n33083_o = n33037_o ? n33082_o : n33067_o;
  assign n33084_o = n33068_o[25:14];
  assign n33085_o = mmcr0[25:14];
  /* pmu.vhdl:156:17  */
  assign n33086_o = n33037_o ? n33084_o : n33085_o;
  assign n33087_o = n33068_o[26];
  /* pmu.vhdl:156:17  */
  assign n33088_o = n33037_o ? n33087_o : n33052_o;
  assign n33089_o = n33068_o[30:27];
  assign n33090_o = mmcr0[30:27];
  /* pmu.vhdl:156:17  */
  assign n33091_o = n33037_o ? n33089_o : n33090_o;
  assign n33092_o = n33068_o[31];
  /* pmu.vhdl:156:17  */
  assign n33093_o = n33037_o ? n33092_o : n33060_o;
  /* pmu.vhdl:173:25  */
  assign n33094_o = n32886_o[1];
  /* pmu.vhdl:173:53  */
  assign n33095_o = n32886_o[5:2];
  /* pmu.vhdl:173:66  */
  assign n33097_o = n33095_o == 4'b1110;
  /* pmu.vhdl:173:37  */
  assign n33098_o = n33094_o & n33097_o;
  /* pmu.vhdl:174:35  */
  assign n33099_o = n32886_o[70:7];
  /* pmu.vhdl:173:17  */
  assign n33100_o = n33098_o ? n33099_o : mmcr1;
  /* pmu.vhdl:176:25  */
  assign n33101_o = n32886_o[1];
  /* pmu.vhdl:176:53  */
  assign n33102_o = n32886_o[5:2];
  /* pmu.vhdl:176:66  */
  assign n33104_o = n33102_o == 4'b0001;
  /* pmu.vhdl:176:37  */
  assign n33105_o = n33101_o & n33104_o;
  /* pmu.vhdl:177:35  */
  assign n33106_o = n32886_o[70:7];
  /* pmu.vhdl:176:17  */
  assign n33107_o = n33105_o ? n33106_o : mmcr2;
  /* pmu.vhdl:179:25  */
  assign n33108_o = n32886_o[1];
  /* pmu.vhdl:179:53  */
  assign n33109_o = n32886_o[5:2];
  /* pmu.vhdl:179:66  */
  assign n33111_o = n33109_o == 4'b0010;
  /* pmu.vhdl:179:37  */
  assign n33112_o = n33108_o & n33111_o;
  assign n33115_o = n32886_o[70:8];
  assign n33116_o = {n33115_o, 1'b0};
  /* pmu.vhdl:179:17  */
  assign n33117_o = n33112_o ? n33116_o : mmcra;
  /* pmu.vhdl:184:25  */
  assign n33118_o = n32886_o[1];
  /* pmu.vhdl:184:53  */
  assign n33119_o = n32886_o[5:2];
  /* pmu.vhdl:184:66  */
  assign n33121_o = n33119_o == 4'b1100;
  /* pmu.vhdl:184:37  */
  assign n33122_o = n33118_o & n33121_o;
  /* pmu.vhdl:185:34  */
  assign n33123_o = n32886_o[70:7];
  /* pmu.vhdl:187:34  */
  assign n33124_o = n32886_o[141:78];
  /* pmu.vhdl:186:17  */
  assign n33125_o = doalert ? n33124_o : siar;
  /* pmu.vhdl:184:17  */
  assign n33126_o = n33122_o ? n33123_o : n33125_o;
  /* pmu.vhdl:189:25  */
  assign n33127_o = n32886_o[1];
  /* pmu.vhdl:189:53  */
  assign n33128_o = n32886_o[5:2];
  /* pmu.vhdl:189:66  */
  assign n33130_o = n33128_o == 4'b1101;
  /* pmu.vhdl:189:37  */
  assign n33131_o = n33127_o & n33130_o;
  /* pmu.vhdl:190:34  */
  assign n33132_o = n32886_o[70:7];
  /* pmu.vhdl:192:34  */
  assign n33133_o = n32886_o[205:142];
  /* pmu.vhdl:191:17  */
  assign n33134_o = doalert ? n33133_o : sdar;
  /* pmu.vhdl:189:17  */
  assign n33135_o = n33131_o ? n33132_o : n33134_o;
  /* pmu.vhdl:194:25  */
  assign n33136_o = n32886_o[1];
  /* pmu.vhdl:194:53  */
  assign n33137_o = n32886_o[5:2];
  /* pmu.vhdl:194:66  */
  assign n33139_o = n33137_o == 4'b0000;
  /* pmu.vhdl:194:37  */
  assign n33140_o = n33136_o & n33139_o;
  /* pmu.vhdl:195:34  */
  assign n33141_o = n32886_o[70:7];
  /* pmu.vhdl:198:47  */
  assign n33142_o = n32886_o[76];
  assign n33144_o = n33143_o[63:26];
  assign n33147_o = n33143_o[24:23];
  /* pmu.vhdl:200:46  */
  assign n33149_o = n32886_o[206];
  assign n33150_o = n33143_o[20:0];
  assign n33151_o = {n33144_o, n33142_o, n33147_o, 1'b1, n33149_o, n33150_o};
  /* pmu.vhdl:196:17  */
  assign n33152_o = doalert ? n33151_o : sier;
  /* pmu.vhdl:194:17  */
  assign n33153_o = n33140_o ? n33141_o : n33152_o;
  assign n33154_o = {n32957_o, n32972_o, n32987_o, n33002_o, n33017_o, n33032_o};
  /* pmu.vhdl:146:13  */
  assign n33155_o = rst ? pmcs : n33154_o;
  assign n33156_o = {n33093_o, n33091_o, n33088_o, n33086_o, n33083_o, n33081_o, n33078_o, n33076_o, n33073_o, n33071_o};
  /* pmu.vhdl:146:13  */
  assign n33158_o = rst ? 32'b10000000000000000000000000000000 : n33156_o;
  /* pmu.vhdl:146:13  */
  assign n33159_o = rst ? mmcr1 : n33100_o;
  /* pmu.vhdl:146:13  */
  assign n33160_o = rst ? mmcr2 : n33107_o;
  /* pmu.vhdl:146:13  */
  assign n33161_o = rst ? mmcra : n33117_o;
  /* pmu.vhdl:146:13  */
  assign n33162_o = rst ? siar : n33126_o;
  /* pmu.vhdl:146:13  */
  assign n33163_o = rst ? sdar : n33135_o;
  /* pmu.vhdl:146:13  */
  assign n33164_o = rst ? sier : n33153_o;
  /* pmu.vhdl:203:29  */
  assign n33165_o = n32886_o[74:71];
  /* pmu.vhdl:219:24  */
  assign n33184_o = n32886_o[74:71];
  /* pmu.vhdl:219:35  */
  assign n33185_o = ~prev_tb;
  /* pmu.vhdl:219:31  */
  assign n33186_o = n33184_o & n33185_o;
  /* pmu.vhdl:220:54  */
  assign n33187_o = mmcr0[24:23];
  /* pmu.vhdl:220:29  */
  assign n33188_o = {29'b0, n33187_o};  //  uext
  /* pmu.vhdl:220:27  */
  assign n33189_o = {1'b0, n33188_o};  //  uext
  /* pmu.vhdl:220:27  */
  assign n33191_o = 32'b00000000000000000000000000000011 - n33189_o;
  /* pmu.vhdl:220:27  */
  assign n33192_o = n33191_o[1:0];  // trunc
  /* pmu.vhdl:221:33  */
  assign n33195_o = mmcr0[22];
  /* pmu.vhdl:221:24  */
  assign n33196_o = n33602_o & n33195_o;
  /* pmu.vhdl:221:9  */
  assign n33199_o = n33196_o ? 1'b1 : 1'b0;
  /* pmu.vhdl:226:17  */
  assign n33201_o = mmcr0[15];
  /* pmu.vhdl:226:49  */
  assign n33202_o = pmcs[191];
  /* pmu.vhdl:226:38  */
  assign n33203_o = n33201_o & n33202_o;
  /* pmu.vhdl:226:9  */
  assign n33205_o = n33203_o ? 1'b1 : n33199_o;
  /* pmu.vhdl:229:17  */
  assign n33206_o = mmcr0[14];
  /* pmu.vhdl:230:21  */
  assign n33207_o = pmcs[159];
  /* pmu.vhdl:230:36  */
  assign n33208_o = pmcs[127];
  /* pmu.vhdl:230:26  */
  assign n33209_o = n33207_o | n33208_o;
  /* pmu.vhdl:230:51  */
  assign n33210_o = pmcs[95];
  /* pmu.vhdl:230:41  */
  assign n33211_o = n33209_o | n33210_o;
  /* pmu.vhdl:229:38  */
  assign n33212_o = n33206_o & n33211_o;
  /* pmu.vhdl:229:9  */
  assign n33214_o = n33212_o ? 1'b1 : n33205_o;
  /* pmu.vhdl:233:17  */
  assign n33215_o = mmcr0[14];
  /* pmu.vhdl:234:18  */
  assign n33216_o = mmcr0[19:18];
  /* pmu.vhdl:234:53  */
  assign n33218_o = n33216_o != 2'b11;
  /* pmu.vhdl:233:38  */
  assign n33219_o = n33215_o & n33218_o;
  /* pmu.vhdl:235:21  */
  assign n33220_o = pmcs[63];
  /* pmu.vhdl:235:36  */
  assign n33221_o = pmcs[31];
  /* pmu.vhdl:235:26  */
  assign n33222_o = n33220_o | n33221_o;
  /* pmu.vhdl:234:61  */
  assign n33223_o = n33219_o & n33222_o;
  /* pmu.vhdl:233:9  */
  assign n33225_o = n33223_o ? 1'b1 : n33214_o;
  /* pmu.vhdl:242:19  */
  assign n33226_o = mmcr1[31:24];
  /* pmu.vhdl:243:13  */
  assign n33229_o = n33226_o == 8'b11110000;
  /* pmu.vhdl:247:32  */
  assign n33230_o = n32886_o[227:207];
  /* pmu.vhdl:247:38  */
  assign n33231_o = n33230_o[3];
  /* pmu.vhdl:246:13  */
  assign n33233_o = n33226_o == 8'b11110010;
  /* pmu.vhdl:246:24  */
  assign n33235_o = n33226_o == 8'b11111110;
  /* pmu.vhdl:246:24  */
  assign n33236_o = n33233_o | n33235_o;
  /* pmu.vhdl:249:32  */
  assign n33237_o = n32886_o[227:207];
  /* pmu.vhdl:249:38  */
  assign n33238_o = n33237_o[4];
  /* pmu.vhdl:248:13  */
  assign n33240_o = n33226_o == 8'b11110100;
  /* pmu.vhdl:251:32  */
  assign n33241_o = n32886_o[227:207];
  /* pmu.vhdl:251:38  */
  assign n33242_o = n33241_o[10];
  /* pmu.vhdl:250:13  */
  assign n33244_o = n33226_o == 8'b11110110;
  /* pmu.vhdl:253:32  */
  assign n33245_o = n32886_o[227:207];
  /* pmu.vhdl:253:38  */
  assign n33246_o = n33245_o[0];
  /* pmu.vhdl:252:13  */
  assign n33248_o = n33226_o == 8'b11111000;
  /* pmu.vhdl:255:32  */
  assign n33249_o = n32886_o[77];
  /* pmu.vhdl:254:13  */
  assign n33251_o = n33226_o == 8'b11111010;
  /* pmu.vhdl:257:32  */
  assign n33252_o = n32886_o[227:207];
  /* pmu.vhdl:257:38  */
  assign n33253_o = n33252_o[5];
  /* pmu.vhdl:256:13  */
  assign n33255_o = n33226_o == 8'b11111100;
  assign n33256_o = {n33255_o, n33251_o, n33248_o, n33244_o, n33240_o, n33236_o, n33229_o};
  /* pmu.vhdl:242:9  */
  always @*
    case (n33256_o)
      7'b1000000: n33258_o = n33253_o;
      7'b0100000: n33258_o = n33249_o;
      7'b0010000: n33258_o = n33246_o;
      7'b0001000: n33258_o = n33242_o;
      7'b0000100: n33258_o = n33238_o;
      7'b0000010: n33258_o = n33231_o;
      7'b0000001: n33258_o = 1'b1;
      default: n33258_o = 1'b0;
    endcase
  /* pmu.vhdl:242:9  */
  always @*
    case (n33256_o)
      7'b1000000: n33263_o = 1'b0;
      7'b0100000: n33263_o = 1'b0;
      7'b0010000: n33263_o = 1'b0;
      7'b0001000: n33263_o = 1'b0;
      7'b0000100: n33263_o = 1'b0;
      7'b0000010: n33263_o = 1'b0;
      7'b0000001: n33263_o = 1'b1;
      default: n33263_o = 1'b0;
    endcase
  /* pmu.vhdl:261:19  */
  assign n33265_o = mmcr1[23:16];
  /* pmu.vhdl:263:32  */
  assign n33266_o = n32886_o[227:207];
  /* pmu.vhdl:263:38  */
  assign n33267_o = n33266_o[6];
  /* pmu.vhdl:262:13  */
  assign n33269_o = n33265_o == 8'b11110000;
  /* pmu.vhdl:265:32  */
  assign n33270_o = n32886_o[227:207];
  /* pmu.vhdl:265:38  */
  assign n33271_o = n33270_o[1];
  /* pmu.vhdl:264:13  */
  assign n33273_o = n33265_o == 8'b11110010;
  /* pmu.vhdl:267:32  */
  assign n33274_o = n32886_o[77];
  /* pmu.vhdl:266:13  */
  assign n33276_o = n33265_o == 8'b11110100;
  /* pmu.vhdl:269:32  */
  assign n33277_o = n32886_o[227:207];
  /* pmu.vhdl:269:38  */
  assign n33278_o = n33277_o[18];
  /* pmu.vhdl:268:13  */
  assign n33280_o = n33265_o == 8'b11110110;
  /* pmu.vhdl:271:32  */
  assign n33281_o = n32886_o[227:207];
  /* pmu.vhdl:271:38  */
  assign n33282_o = n33281_o[2];
  /* pmu.vhdl:270:13  */
  assign n33284_o = n33265_o == 8'b11111000;
  /* pmu.vhdl:273:32  */
  assign n33285_o = n32886_o[227:207];
  /* pmu.vhdl:273:38  */
  assign n33286_o = n33285_o[7];
  /* pmu.vhdl:272:13  */
  assign n33288_o = n33265_o == 8'b11111010;
  /* pmu.vhdl:275:32  */
  assign n33289_o = n32886_o[227:207];
  /* pmu.vhdl:275:38  */
  assign n33290_o = n33289_o[12];
  /* pmu.vhdl:274:13  */
  assign n33292_o = n33265_o == 8'b11111100;
  /* pmu.vhdl:277:32  */
  assign n33293_o = n32886_o[227:207];
  /* pmu.vhdl:277:38  */
  assign n33294_o = n33293_o[13];
  /* pmu.vhdl:276:13  */
  assign n33296_o = n33265_o == 8'b11111110;
  assign n33297_o = {n33296_o, n33292_o, n33288_o, n33284_o, n33280_o, n33276_o, n33273_o, n33269_o};
  assign n33298_o = n33259_o[4];
  /* pmu.vhdl:261:9  */
  always @*
    case (n33297_o)
      8'b10000000: n33299_o = n33294_o;
      8'b01000000: n33299_o = n33290_o;
      8'b00100000: n33299_o = n33286_o;
      8'b00010000: n33299_o = n33282_o;
      8'b00001000: n33299_o = n33278_o;
      8'b00000100: n33299_o = n33274_o;
      8'b00000010: n33299_o = n33271_o;
      8'b00000001: n33299_o = n33267_o;
      default: n33299_o = n33298_o;
    endcase
  /* pmu.vhdl:281:19  */
  assign n33301_o = mmcr1[15:8];
  /* pmu.vhdl:283:32  */
  assign n33302_o = n32886_o[227:207];
  /* pmu.vhdl:283:38  */
  assign n33303_o = n33302_o[16];
  /* pmu.vhdl:282:13  */
  assign n33305_o = n33301_o == 8'b11110000;
  /* pmu.vhdl:285:32  */
  assign n33306_o = n32886_o[227:207];
  /* pmu.vhdl:285:38  */
  assign n33307_o = n33306_o[1];
  /* pmu.vhdl:284:13  */
  assign n33309_o = n33301_o == 8'b11110010;
  /* pmu.vhdl:287:32  */
  assign n33310_o = n32886_o[227:207];
  /* pmu.vhdl:287:38  */
  assign n33311_o = n33310_o[3];
  /* pmu.vhdl:287:62  */
  assign n33312_o = n32886_o[77];
  /* pmu.vhdl:287:53  */
  assign n33313_o = n33311_o & n33312_o;
  /* pmu.vhdl:286:13  */
  assign n33315_o = n33301_o == 8'b11110100;
  /* pmu.vhdl:289:32  */
  assign n33316_o = n32886_o[227:207];
  /* pmu.vhdl:289:38  */
  assign n33317_o = n33316_o[15];
  /* pmu.vhdl:288:13  */
  assign n33319_o = n33301_o == 8'b11110110;
  /* pmu.vhdl:290:13  */
  assign n33321_o = n33301_o == 8'b11111000;
  /* pmu.vhdl:293:32  */
  assign n33322_o = n32886_o[227:207];
  /* pmu.vhdl:293:38  */
  assign n33323_o = n33322_o[17];
  /* pmu.vhdl:292:13  */
  assign n33325_o = n33301_o == 8'b11111110;
  assign n33326_o = {n33325_o, n33321_o, n33319_o, n33315_o, n33309_o, n33305_o};
  assign n33327_o = n33259_o[3];
  /* pmu.vhdl:281:9  */
  always @*
    case (n33326_o)
      6'b100000: n33328_o = n33323_o;
      6'b010000: n33328_o = n33602_o;
      6'b001000: n33328_o = n33317_o;
      6'b000100: n33328_o = n33313_o;
      6'b000010: n33328_o = n33307_o;
      6'b000001: n33328_o = n33303_o;
      default: n33328_o = n33327_o;
    endcase
  /* pmu.vhdl:297:19  */
  assign n33330_o = mmcr1[7:0];
  /* pmu.vhdl:299:32  */
  assign n33331_o = n32886_o[227:207];
  /* pmu.vhdl:299:38  */
  assign n33332_o = n33331_o[14];
  /* pmu.vhdl:298:13  */
  assign n33334_o = n33330_o == 8'b11110000;
  /* pmu.vhdl:301:32  */
  assign n33335_o = n32886_o[227:207];
  /* pmu.vhdl:301:38  */
  assign n33336_o = n33335_o[1];
  /* pmu.vhdl:300:13  */
  assign n33338_o = n33330_o == 8'b11110010;
  /* pmu.vhdl:303:32  */
  assign n33339_o = n32886_o[77];
  /* pmu.vhdl:302:13  */
  assign n33341_o = n33330_o == 8'b11110100;
  /* pmu.vhdl:305:32  */
  assign n33342_o = n32886_o[227:207];
  /* pmu.vhdl:305:38  */
  assign n33343_o = n33342_o[8];
  /* pmu.vhdl:304:13  */
  assign n33345_o = n33330_o == 8'b11110110;
  /* pmu.vhdl:307:32  */
  assign n33346_o = n32886_o[227:207];
  /* pmu.vhdl:307:38  */
  assign n33347_o = n33346_o[9];
  /* pmu.vhdl:306:13  */
  assign n33349_o = n33330_o == 8'b11111000;
  /* pmu.vhdl:309:32  */
  assign n33350_o = n32886_o[227:207];
  /* pmu.vhdl:309:38  */
  assign n33351_o = n33350_o[3];
  /* pmu.vhdl:309:62  */
  assign n33352_o = n32886_o[77];
  /* pmu.vhdl:309:53  */
  assign n33353_o = n33351_o & n33352_o;
  /* pmu.vhdl:308:13  */
  assign n33355_o = n33330_o == 8'b11111010;
  /* pmu.vhdl:311:32  */
  assign n33356_o = n32886_o[227:207];
  /* pmu.vhdl:311:38  */
  assign n33357_o = n33356_o[11];
  /* pmu.vhdl:310:13  */
  assign n33359_o = n33330_o == 8'b11111100;
  /* pmu.vhdl:313:32  */
  assign n33360_o = n32886_o[227:207];
  /* pmu.vhdl:313:38  */
  assign n33361_o = n33360_o[19];
  /* pmu.vhdl:312:13  */
  assign n33363_o = n33330_o == 8'b11111110;
  assign n33364_o = {n33363_o, n33359_o, n33355_o, n33349_o, n33345_o, n33341_o, n33338_o, n33334_o};
  assign n33365_o = n33259_o[2];
  /* pmu.vhdl:297:9  */
  always @*
    case (n33364_o)
      8'b10000000: n33366_o = n33361_o;
      8'b01000000: n33366_o = n33357_o;
      8'b00100000: n33366_o = n33353_o;
      8'b00010000: n33366_o = n33347_o;
      8'b00001000: n33366_o = n33343_o;
      8'b00000100: n33366_o = n33339_o;
      8'b00000010: n33366_o = n33336_o;
      8'b00000001: n33366_o = n33332_o;
      default: n33366_o = n33365_o;
    endcase
  /* pmu.vhdl:317:25  */
  assign n33368_o = mmcr0[8];
  /* pmu.vhdl:317:49  */
  assign n33369_o = n32886_o[77];
  /* pmu.vhdl:317:41  */
  assign n33370_o = n33368_o | n33369_o;
  /* pmu.vhdl:317:63  */
  assign n33371_o = n32886_o[227:207];
  /* pmu.vhdl:317:69  */
  assign n33372_o = n33371_o[3];
  /* pmu.vhdl:317:54  */
  assign n33373_o = n33370_o & n33372_o;
  /* pmu.vhdl:318:24  */
  assign n33375_o = mmcr0[8];
  /* pmu.vhdl:318:48  */
  assign n33376_o = n32886_o[77];
  /* pmu.vhdl:318:40  */
  assign n33377_o = n33375_o | n33376_o;
  /* pmu.vhdl:321:24  */
  assign n33378_o = mmcr0[31];
  /* pmu.vhdl:322:25  */
  assign n33379_o = mmcr0[30];
  /* pmu.vhdl:322:50  */
  assign n33380_o = n32886_o[76];
  /* pmu.vhdl:322:41  */
  assign n33381_o = ~n33380_o;
  /* pmu.vhdl:322:37  */
  assign n33382_o = n33379_o & n33381_o;
  /* pmu.vhdl:321:35  */
  assign n33383_o = n33378_o | n33382_o;
  /* pmu.vhdl:323:25  */
  assign n33384_o = mmcr0[29];
  /* pmu.vhdl:323:50  */
  assign n33385_o = mmcr0[12];
  /* pmu.vhdl:323:41  */
  assign n33386_o = ~n33385_o;
  /* pmu.vhdl:323:37  */
  assign n33387_o = n33384_o & n33386_o;
  /* pmu.vhdl:323:72  */
  assign n33388_o = n32886_o[76];
  /* pmu.vhdl:323:63  */
  assign n33389_o = n33387_o & n33388_o;
  /* pmu.vhdl:322:58  */
  assign n33390_o = n33383_o | n33389_o;
  /* pmu.vhdl:324:29  */
  assign n33391_o = mmcr0[29];
  /* pmu.vhdl:324:20  */
  assign n33392_o = ~n33391_o;
  /* pmu.vhdl:324:50  */
  assign n33393_o = mmcr0[12];
  /* pmu.vhdl:324:41  */
  assign n33394_o = n33392_o & n33393_o;
  /* pmu.vhdl:324:72  */
  assign n33395_o = n32886_o[76];
  /* pmu.vhdl:324:63  */
  assign n33396_o = n33394_o & n33395_o;
  /* pmu.vhdl:323:80  */
  assign n33397_o = n33390_o | n33396_o;
  /* pmu.vhdl:325:25  */
  assign n33398_o = mmcr0[28];
  /* pmu.vhdl:325:47  */
  assign n33399_o = n32886_o[75];
  /* pmu.vhdl:325:38  */
  assign n33400_o = n33398_o & n33399_o;
  /* pmu.vhdl:324:80  */
  assign n33401_o = n33397_o | n33400_o;
  /* pmu.vhdl:326:25  */
  assign n33402_o = mmcr0[27];
  /* pmu.vhdl:326:51  */
  assign n33403_o = n32886_o[75];
  /* pmu.vhdl:326:42  */
  assign n33404_o = ~n33403_o;
  /* pmu.vhdl:326:38  */
  assign n33405_o = n33402_o & n33404_o;
  /* pmu.vhdl:325:56  */
  assign n33406_o = n33401_o | n33405_o;
  /* pmu.vhdl:328:33  */
  assign n33407_o = mmcr0[5];
  /* pmu.vhdl:328:25  */
  assign n33408_o = n33406_o | n33407_o;
  /* pmu.vhdl:329:19  */
  assign n33409_o = mmcr0[1];
  /* pmu.vhdl:329:49  */
  assign n33410_o = n32886_o[77];
  /* pmu.vhdl:329:53  */
  assign n33411_o = ~n33410_o;
  /* pmu.vhdl:329:40  */
  assign n33412_o = n33409_o & n33411_o;
  /* pmu.vhdl:329:70  */
  assign n33413_o = ~n33263_o;
  /* pmu.vhdl:329:59  */
  assign n33414_o = n33412_o & n33413_o;
  /* pmu.vhdl:328:53  */
  assign n33415_o = n33408_o | n33414_o;
  /* pmu.vhdl:328:9  */
  assign n33417_o = n33415_o ? 1'b0 : n33258_o;
  /* pmu.vhdl:332:33  */
  assign n33418_o = mmcr0[5];
  /* pmu.vhdl:332:25  */
  assign n33419_o = n33406_o | n33418_o;
  /* pmu.vhdl:333:19  */
  assign n33420_o = mmcr0[1];
  /* pmu.vhdl:333:49  */
  assign n33421_o = n32886_o[77];
  /* pmu.vhdl:333:53  */
  assign n33422_o = ~n33421_o;
  /* pmu.vhdl:333:40  */
  assign n33423_o = n33420_o & n33422_o;
  /* pmu.vhdl:332:53  */
  assign n33424_o = n33419_o | n33423_o;
  assign n33426_o = {n33299_o, n33328_o, n33366_o};
  /* pmu.vhdl:332:9  */
  assign n33427_o = n33424_o ? 3'b000 : n33426_o;
  /* pmu.vhdl:336:33  */
  assign n33428_o = mmcr0[4];
  /* pmu.vhdl:336:25  */
  assign n33429_o = n33406_o | n33428_o;
  assign n33431_o = {n33373_o, n33377_o};
  /* pmu.vhdl:336:9  */
  assign n33432_o = n33429_o ? 2'b00 : n33431_o;
  /* pmu.vhdl:339:17  */
  assign n33433_o = mmcr0[13];
  assign n33435_o = {n33427_o, n33432_o};
  /* pmu.vhdl:344:22  */
  assign n33437_o = mmcr2[63];
  /* pmu.vhdl:344:54  */
  assign n33438_o = n32886_o[76];
  /* pmu.vhdl:344:61  */
  assign n33439_o = ~n33438_o;
  /* pmu.vhdl:344:45  */
  assign n33440_o = n33437_o & n33439_o;
  /* pmu.vhdl:345:23  */
  assign n33441_o = mmcr2[62];
  /* pmu.vhdl:345:56  */
  assign n33442_o = n32886_o[76];
  /* pmu.vhdl:345:47  */
  assign n33443_o = n33441_o & n33442_o;
  /* pmu.vhdl:344:68  */
  assign n33444_o = n33440_o | n33443_o;
  /* pmu.vhdl:346:23  */
  assign n33445_o = mmcr2[60];
  /* pmu.vhdl:346:56  */
  assign n33446_o = n32886_o[75];
  /* pmu.vhdl:346:47  */
  assign n33447_o = n33445_o & n33446_o;
  /* pmu.vhdl:345:70  */
  assign n33448_o = n33444_o | n33447_o;
  /* pmu.vhdl:347:23  */
  assign n33449_o = mmcr2[60];
  /* pmu.vhdl:347:56  */
  assign n33450_o = n32886_o[75];
  /* pmu.vhdl:347:47  */
  assign n33451_o = n33449_o & n33450_o;
  /* pmu.vhdl:346:71  */
  assign n33452_o = n33448_o | n33451_o;
  /* pmu.vhdl:344:13  */
  assign n33454_o = n33452_o ? 1'b0 : n33417_o;
  /* pmu.vhdl:344:22  */
  assign n33455_o = mmcr2[54];
  /* pmu.vhdl:344:54  */
  assign n33456_o = n32886_o[76];
  /* pmu.vhdl:344:61  */
  assign n33457_o = ~n33456_o;
  /* pmu.vhdl:344:45  */
  assign n33458_o = n33455_o & n33457_o;
  /* pmu.vhdl:345:23  */
  assign n33459_o = mmcr2[53];
  /* pmu.vhdl:345:56  */
  assign n33460_o = n32886_o[76];
  /* pmu.vhdl:345:47  */
  assign n33461_o = n33459_o & n33460_o;
  /* pmu.vhdl:344:68  */
  assign n33462_o = n33458_o | n33461_o;
  /* pmu.vhdl:346:23  */
  assign n33463_o = mmcr2[51];
  /* pmu.vhdl:346:56  */
  assign n33464_o = n32886_o[75];
  /* pmu.vhdl:346:47  */
  assign n33465_o = n33463_o & n33464_o;
  /* pmu.vhdl:345:70  */
  assign n33466_o = n33462_o | n33465_o;
  /* pmu.vhdl:347:23  */
  assign n33467_o = mmcr2[51];
  /* pmu.vhdl:347:56  */
  assign n33468_o = n32886_o[75];
  /* pmu.vhdl:347:47  */
  assign n33469_o = n33467_o & n33468_o;
  /* pmu.vhdl:346:71  */
  assign n33470_o = n33466_o | n33469_o;
  assign n33472_o = n33434_o[4];
  assign n33473_o = n33435_o[4];
  /* pmu.vhdl:339:9  */
  assign n33474_o = n33433_o ? n33472_o : n33473_o;
  /* pmu.vhdl:344:13  */
  assign n33475_o = n33470_o ? 1'b0 : n33474_o;
  /* pmu.vhdl:344:22  */
  assign n33479_o = mmcr2[45];
  /* pmu.vhdl:344:54  */
  assign n33480_o = n32886_o[76];
  /* pmu.vhdl:344:61  */
  assign n33481_o = ~n33480_o;
  /* pmu.vhdl:344:45  */
  assign n33482_o = n33479_o & n33481_o;
  /* pmu.vhdl:345:23  */
  assign n33483_o = mmcr2[44];
  /* pmu.vhdl:345:56  */
  assign n33484_o = n32886_o[76];
  /* pmu.vhdl:345:47  */
  assign n33485_o = n33483_o & n33484_o;
  /* pmu.vhdl:344:68  */
  assign n33486_o = n33482_o | n33485_o;
  /* pmu.vhdl:346:23  */
  assign n33487_o = mmcr2[42];
  /* pmu.vhdl:346:56  */
  assign n33488_o = n32886_o[75];
  /* pmu.vhdl:346:47  */
  assign n33489_o = n33487_o & n33488_o;
  /* pmu.vhdl:345:70  */
  assign n33490_o = n33486_o | n33489_o;
  /* pmu.vhdl:347:23  */
  assign n33491_o = mmcr2[42];
  /* pmu.vhdl:347:56  */
  assign n33492_o = n32886_o[75];
  /* pmu.vhdl:347:47  */
  assign n33493_o = n33491_o & n33492_o;
  /* pmu.vhdl:346:71  */
  assign n33494_o = n33490_o | n33493_o;
  assign n33496_o = n33434_o[3];
  assign n33497_o = n33435_o[3];
  /* pmu.vhdl:339:9  */
  assign n33498_o = n33433_o ? n33496_o : n33497_o;
  /* pmu.vhdl:344:13  */
  assign n33499_o = n33494_o ? 1'b0 : n33498_o;
  /* pmu.vhdl:344:22  */
  assign n33503_o = mmcr2[36];
  /* pmu.vhdl:344:54  */
  assign n33504_o = n32886_o[76];
  /* pmu.vhdl:344:61  */
  assign n33505_o = ~n33504_o;
  /* pmu.vhdl:344:45  */
  assign n33506_o = n33503_o & n33505_o;
  /* pmu.vhdl:345:23  */
  assign n33507_o = mmcr2[35];
  /* pmu.vhdl:345:56  */
  assign n33508_o = n32886_o[76];
  /* pmu.vhdl:345:47  */
  assign n33509_o = n33507_o & n33508_o;
  /* pmu.vhdl:344:68  */
  assign n33510_o = n33506_o | n33509_o;
  /* pmu.vhdl:346:23  */
  assign n33511_o = mmcr2[33];
  /* pmu.vhdl:346:56  */
  assign n33512_o = n32886_o[75];
  /* pmu.vhdl:346:47  */
  assign n33513_o = n33511_o & n33512_o;
  /* pmu.vhdl:345:70  */
  assign n33514_o = n33510_o | n33513_o;
  /* pmu.vhdl:347:23  */
  assign n33515_o = mmcr2[33];
  /* pmu.vhdl:347:56  */
  assign n33516_o = n32886_o[75];
  /* pmu.vhdl:347:47  */
  assign n33517_o = n33515_o & n33516_o;
  /* pmu.vhdl:346:71  */
  assign n33518_o = n33514_o | n33517_o;
  assign n33520_o = n33434_o[2];
  assign n33521_o = n33435_o[2];
  /* pmu.vhdl:339:9  */
  assign n33522_o = n33433_o ? n33520_o : n33521_o;
  /* pmu.vhdl:344:13  */
  assign n33523_o = n33518_o ? 1'b0 : n33522_o;
  /* pmu.vhdl:344:22  */
  assign n33527_o = mmcr2[27];
  /* pmu.vhdl:344:54  */
  assign n33528_o = n32886_o[76];
  /* pmu.vhdl:344:61  */
  assign n33529_o = ~n33528_o;
  /* pmu.vhdl:344:45  */
  assign n33530_o = n33527_o & n33529_o;
  /* pmu.vhdl:345:23  */
  assign n33531_o = mmcr2[26];
  /* pmu.vhdl:345:56  */
  assign n33532_o = n32886_o[76];
  /* pmu.vhdl:345:47  */
  assign n33533_o = n33531_o & n33532_o;
  /* pmu.vhdl:344:68  */
  assign n33534_o = n33530_o | n33533_o;
  /* pmu.vhdl:346:23  */
  assign n33535_o = mmcr2[24];
  /* pmu.vhdl:346:56  */
  assign n33536_o = n32886_o[75];
  /* pmu.vhdl:346:47  */
  assign n33537_o = n33535_o & n33536_o;
  /* pmu.vhdl:345:70  */
  assign n33538_o = n33534_o | n33537_o;
  /* pmu.vhdl:347:23  */
  assign n33539_o = mmcr2[24];
  /* pmu.vhdl:347:56  */
  assign n33540_o = n32886_o[75];
  /* pmu.vhdl:347:47  */
  assign n33541_o = n33539_o & n33540_o;
  /* pmu.vhdl:346:71  */
  assign n33542_o = n33538_o | n33541_o;
  assign n33544_o = n33434_o[1];
  assign n33545_o = n33435_o[1];
  /* pmu.vhdl:339:9  */
  assign n33546_o = n33433_o ? n33544_o : n33545_o;
  /* pmu.vhdl:344:13  */
  assign n33547_o = n33542_o ? 1'b0 : n33546_o;
  assign n33548_o = n33434_o[0];
  assign n33549_o = n33435_o[0];
  /* pmu.vhdl:339:9  */
  assign n33550_o = n33433_o ? n33548_o : n33549_o;
  /* pmu.vhdl:344:22  */
  assign n33551_o = mmcr2[18];
  /* pmu.vhdl:344:54  */
  assign n33552_o = n32886_o[76];
  /* pmu.vhdl:344:61  */
  assign n33553_o = ~n33552_o;
  /* pmu.vhdl:344:45  */
  assign n33554_o = n33551_o & n33553_o;
  /* pmu.vhdl:345:23  */
  assign n33555_o = mmcr2[17];
  /* pmu.vhdl:345:56  */
  assign n33556_o = n32886_o[76];
  /* pmu.vhdl:345:47  */
  assign n33557_o = n33555_o & n33556_o;
  /* pmu.vhdl:344:68  */
  assign n33558_o = n33554_o | n33557_o;
  /* pmu.vhdl:346:23  */
  assign n33559_o = mmcr2[15];
  /* pmu.vhdl:346:56  */
  assign n33560_o = n32886_o[75];
  /* pmu.vhdl:346:47  */
  assign n33561_o = n33559_o & n33560_o;
  /* pmu.vhdl:345:70  */
  assign n33562_o = n33558_o | n33561_o;
  /* pmu.vhdl:347:23  */
  assign n33563_o = mmcr2[15];
  /* pmu.vhdl:347:56  */
  assign n33564_o = n32886_o[75];
  /* pmu.vhdl:347:47  */
  assign n33565_o = n33563_o & n33564_o;
  /* pmu.vhdl:346:71  */
  assign n33566_o = n33562_o | n33565_o;
  /* pmu.vhdl:344:13  */
  assign n33568_o = n33566_o ? 1'b0 : n33550_o;
  /* pmu.vhdl:355:17  */
  assign n33569_o = mmcr0[19:18];
  /* pmu.vhdl:355:52  */
  assign n33571_o = n33569_o == 2'b11;
  /* pmu.vhdl:356:28  */
  assign n33572_o = n32886_o[77];
  /* pmu.vhdl:356:41  */
  assign n33573_o = n32886_o[227:207];
  /* pmu.vhdl:356:47  */
  assign n33574_o = n33573_o[3];
  /* pmu.vhdl:356:32  */
  assign n33575_o = n33572_o & n33574_o;
  /* pmu.vhdl:357:28  */
  assign n33576_o = n32886_o[77];
  assign n33577_o = {n33575_o, n33576_o};
  assign n33578_o = {n33547_o, n33568_o};
  /* pmu.vhdl:355:9  */
  assign n33579_o = n33571_o ? n33577_o : n33578_o;
  assign n33580_o = {n33454_o, n33475_o, n33499_o, n33523_o, n33579_o};
  /* pmu.vhdl:362:35  */
  assign n33581_o = mmcr0[26];
  /* pmu.vhdl:362:26  */
  assign n33582_o = n33225_o & n33581_o;
  /* pmu.vhdl:145:9  */
  always @(posedge clk)
    n33587_q <= n33155_o;
  /* pmu.vhdl:145:9  */
  always @(posedge clk)
    n33588_q <= n33158_o;
  /* pmu.vhdl:145:9  */
  always @(posedge clk)
    n33589_q <= n33159_o;
  /* pmu.vhdl:145:9  */
  always @(posedge clk)
    n33590_q <= n33160_o;
  /* pmu.vhdl:145:9  */
  always @(posedge clk)
    n33591_q <= n33161_o;
  /* pmu.vhdl:145:9  */
  always @(posedge clk)
    n33592_q <= n33162_o;
  /* pmu.vhdl:145:9  */
  always @(posedge clk)
    n33593_q <= n33163_o;
  /* pmu.vhdl:145:9  */
  always @(posedge clk)
    n33594_q <= n33164_o;
  /* pmu.vhdl:145:9  */
  always @(posedge clk)
    n33595_q <= n33165_o;
  /* pmu.vhdl:145:9  */
  assign n33596_o = {n32940_o, n32939_o};
  assign n33597_o = n33186_o[0];
  /* pmu.vhdl:14:9  */
  assign n33598_o = n33186_o[1];
  assign n33599_o = n33186_o[2];
  assign n33600_o = n33186_o[3];
  /* pmu.vhdl:220:24  */
  assign n33601_o = n33192_o[1:0];
  /* pmu.vhdl:220:24  */
  always @*
    case (n33601_o)
      2'b00: n33602_o = n33597_o;
      2'b01: n33602_o = n33598_o;
      2'b10: n33602_o = n33599_o;
      2'b11: n33602_o = n33600_o;
    endcase
endmodule

module random
  (input  clk,
   output [63:0] data,
   output [63:0] raw,
   output err);
  localparam [63:0] n32883_o = 64'b1111111111111111111111111111111111111111111111111111111111111111;
  localparam [63:0] n32884_o = 64'b1111111111111111111111111111111111111111111111111111111111111111;
  localparam n32885_o = 1'b1;
  assign data = n32883_o;
  assign raw = n32884_o;
  assign err = n32885_o;
endmodule

module divider
  (input  clk,
   input  rst,
   input  d_in_valid,
   input  [63:0] d_in_dividend,
   input  [63:0] d_in_divisor,
   input  d_in_is_signed,
   input  d_in_is_32bit,
   input  d_in_is_extended,
   input  d_in_is_modulus,
   input  d_in_neg_result,
   output d_out_valid,
   output [63:0] d_out_write_reg_data,
   output d_out_overflow);
  wire [133:0] n32686_o;
  wire n32688_o;
  wire [63:0] n32689_o;
  wire n32690_o;
  wire [128:0] dend;
  wire [63:0] div;
  wire [63:0] quot;
  wire [63:0] result;
  wire [64:0] sresult;
  wire [63:0] oresult;
  wire running;
  wire [6:0] count;
  wire neg_result;
  wire is_modulus;
  wire is_32bit;
  wire is_signed;
  wire overflow;
  wire ovf32;
  wire did_ovf;
  wire n32693_o;
  wire n32694_o;
  wire [63:0] n32695_o;
  wire [64:0] n32697_o;
  wire [128:0] n32699_o;
  wire [63:0] n32700_o;
  wire [128:0] n32702_o;
  wire [128:0] n32703_o;
  wire [63:0] n32704_o;
  wire n32705_o;
  wire n32706_o;
  wire n32708_o;
  wire n32709_o;
  wire n32711_o;
  wire n32713_o;
  wire n32714_o;
  wire n32715_o;
  wire [63:0] n32716_o;
  wire n32717_o;
  wire n32718_o;
  wire n32719_o;
  wire n32720_o;
  wire [63:0] n32721_o;
  wire [63:0] n32722_o;
  wire [63:0] n32723_o;
  wire [127:0] n32724_o;
  wire [128:0] n32726_o;
  wire [62:0] n32727_o;
  wire [63:0] n32729_o;
  wire [6:0] n32731_o;
  wire [71:0] n32732_o;
  wire n32734_o;
  wire [3:0] n32735_o;
  wire n32737_o;
  wire n32738_o;
  wire [7:0] n32739_o;
  wire [8:0] n32740_o;
  wire n32741_o;
  wire [120:0] n32742_o;
  wire [128:0] n32744_o;
  wire [55:0] n32745_o;
  wire [63:0] n32747_o;
  wire [6:0] n32749_o;
  wire n32750_o;
  wire n32751_o;
  wire [127:0] n32752_o;
  wire [128:0] n32754_o;
  wire [62:0] n32755_o;
  wire [63:0] n32757_o;
  wire [6:0] n32759_o;
  wire [128:0] n32760_o;
  wire [63:0] n32761_o;
  wire [6:0] n32762_o;
  wire n32763_o;
  wire [128:0] n32764_o;
  wire [63:0] n32765_o;
  wire [6:0] n32766_o;
  wire n32767_o;
  wire [128:0] n32768_o;
  wire [63:0] n32769_o;
  wire n32770_o;
  wire [6:0] n32772_o;
  wire n32773_o;
  wire n32774_o;
  wire [128:0] n32775_o;
  wire [63:0] n32776_o;
  wire [63:0] n32778_o;
  wire n32780_o;
  wire [6:0] n32782_o;
  wire n32783_o;
  wire n32784_o;
  wire n32785_o;
  wire n32787_o;
  wire n32789_o;
  wire n32791_o;
  wire [128:0] n32793_o;
  wire [63:0] n32795_o;
  wire [63:0] n32797_o;
  wire n32799_o;
  wire [6:0] n32801_o;
  wire n32802_o;
  wire n32803_o;
  wire n32804_o;
  wire n32806_o;
  wire n32807_o;
  wire n32808_o;
  wire [63:0] n32823_o;
  wire [63:0] n32824_o;
  wire [64:0] n32826_o;
  wire [64:0] n32827_o;
  wire [64:0] n32829_o;
  wire [64:0] n32830_o;
  wire n32831_o;
  wire n32832_o;
  wire n32833_o;
  wire n32834_o;
  wire n32835_o;
  wire n32836_o;
  wire n32837_o;
  wire n32838_o;
  wire n32839_o;
  wire n32840_o;
  wire n32843_o;
  wire n32844_o;
  wire n32845_o;
  wire n32847_o;
  wire n32848_o;
  wire [31:0] n32849_o;
  wire [63:0] n32851_o;
  wire [63:0] n32852_o;
  wire [63:0] n32853_o;
  wire [63:0] n32855_o;
  wire n32861_o;
  wire n32863_o;
  wire [65:0] n32864_o;
  reg [128:0] n32867_q;
  reg [63:0] n32868_q;
  reg [63:0] n32869_q;
  reg n32870_q;
  reg [6:0] n32871_q;
  reg n32872_q;
  reg n32873_q;
  reg n32874_q;
  reg n32876_q;
  reg n32877_q;
  reg n32878_q;
  reg [65:0] n32879_q;
  assign d_out_valid = n32688_o;
  assign d_out_write_reg_data = n32689_o;
  assign d_out_overflow = n32690_o;
  assign n32686_o = {d_in_neg_result, d_in_is_modulus, d_in_is_extended, d_in_is_32bit, d_in_is_signed, d_in_divisor, d_in_dividend, d_in_valid};
  /* asic/multiply.vhdl:16:9  */
  assign n32688_o = n32879_q[0];
  assign n32689_o = n32879_q[64:1];
  assign n32690_o = n32879_q[65];
  /* divider.vhdl:19:12  */
  assign dend = n32867_q; // (signal)
  /* divider.vhdl:20:12  */
  assign div = n32868_q; // (signal)
  /* divider.vhdl:21:12  */
  assign quot = n32869_q; // (signal)
  /* divider.vhdl:22:12  */
  assign result = n32824_o; // (signal)
  /* divider.vhdl:23:12  */
  assign sresult = n32830_o; // (signal)
  /* divider.vhdl:24:12  */
  assign oresult = n32855_o; // (signal)
  /* divider.vhdl:25:12  */
  assign running = n32870_q; // (signal)
  /* divider.vhdl:26:12  */
  assign count = n32871_q; // (signal)
  /* divider.vhdl:27:12  */
  assign neg_result = n32872_q; // (signal)
  /* divider.vhdl:28:12  */
  assign is_modulus = n32873_q; // (signal)
  /* divider.vhdl:29:12  */
  assign is_32bit = n32874_q; // (signal)
  /* divider.vhdl:31:12  */
  assign is_signed = n32876_q; // (signal)
  /* divider.vhdl:32:12  */
  assign overflow = n32877_q; // (signal)
  /* divider.vhdl:33:12  */
  assign ovf32 = n32878_q; // (signal)
  /* divider.vhdl:34:12  */
  assign did_ovf = n32845_o; // (signal)
  /* divider.vhdl:45:24  */
  assign n32693_o = n32686_o[0];
  /* divider.vhdl:46:25  */
  assign n32694_o = n32686_o[131];
  /* divider.vhdl:47:40  */
  assign n32695_o = n32686_o[64:1];
  /* divider.vhdl:47:33  */
  assign n32697_o = {1'b0, n32695_o};
  /* divider.vhdl:47:49  */
  assign n32699_o = {n32697_o, 64'b0000000000000000000000000000000000000000000000000000000000000000};
  /* divider.vhdl:49:62  */
  assign n32700_o = n32686_o[64:1];
  /* divider.vhdl:49:55  */
  assign n32702_o = {65'b00000000000000000000000000000000000000000000000000000000000000000, n32700_o};
  /* divider.vhdl:46:17  */
  assign n32703_o = n32694_o ? n32699_o : n32702_o;
  /* divider.vhdl:51:38  */
  assign n32704_o = n32686_o[128:65];
  /* divider.vhdl:53:36  */
  assign n32705_o = n32686_o[133];
  /* divider.vhdl:54:36  */
  assign n32706_o = n32686_o[132];
  /* divider.vhdl:56:34  */
  assign n32708_o = n32686_o[130];
  /* divider.vhdl:57:35  */
  assign n32709_o = n32686_o[129];
  /* divider.vhdl:63:26  */
  assign n32711_o = count == 7'b0111111;
  /* divider.vhdl:62:13  */
  assign n32713_o = n32770_o ? 1'b0 : running;
  /* divider.vhdl:66:33  */
  assign n32714_o = quot[63];
  /* divider.vhdl:67:24  */
  assign n32715_o = dend[128];
  /* divider.vhdl:67:52  */
  assign n32716_o = dend[127:64];
  /* divider.vhdl:67:69  */
  assign n32717_o = $unsigned(n32716_o) >= $unsigned(div);
  /* divider.vhdl:67:36  */
  assign n32718_o = n32715_o | n32717_o;
  /* divider.vhdl:68:43  */
  assign n32719_o = quot[31];
  /* divider.vhdl:68:36  */
  assign n32720_o = ovf32 | n32719_o;
  /* divider.vhdl:69:60  */
  assign n32721_o = dend[127:64];
  /* divider.vhdl:69:77  */
  assign n32722_o = n32721_o - div;
  /* divider.vhdl:70:33  */
  assign n32723_o = dend[63:0];
  /* divider.vhdl:69:84  */
  assign n32724_o = {n32722_o, n32723_o};
  /* divider.vhdl:70:47  */
  assign n32726_o = {n32724_o, 1'b0};
  /* divider.vhdl:71:33  */
  assign n32727_o = quot[62:0];
  /* divider.vhdl:71:47  */
  assign n32729_o = {n32727_o, 1'b1};
  /* divider.vhdl:72:36  */
  assign n32731_o = count + 7'b0000001;
  /* divider.vhdl:73:27  */
  assign n32732_o = dend[128:57];
  /* divider.vhdl:73:43  */
  assign n32734_o = n32732_o == 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
  /* divider.vhdl:73:76  */
  assign n32735_o = count[6:3];
  /* divider.vhdl:73:89  */
  assign n32737_o = n32735_o != 4'b0111;
  /* divider.vhdl:73:67  */
  assign n32738_o = n32734_o & n32737_o;
  /* divider.vhdl:75:46  */
  assign n32739_o = quot[31:24];
  /* divider.vhdl:75:40  */
  assign n32740_o = {ovf32, n32739_o};
  /* divider.vhdl:75:30  */
  assign n32741_o = |(n32740_o);
  /* divider.vhdl:76:33  */
  assign n32742_o = dend[120:0];
  /* divider.vhdl:76:48  */
  assign n32744_o = {n32742_o, 8'b00000000};
  /* divider.vhdl:77:33  */
  assign n32745_o = quot[55:0];
  /* divider.vhdl:77:47  */
  assign n32747_o = {n32745_o, 8'b00000000};
  /* divider.vhdl:78:36  */
  assign n32749_o = count + 7'b0001000;
  /* divider.vhdl:80:43  */
  assign n32750_o = quot[31];
  /* divider.vhdl:80:36  */
  assign n32751_o = ovf32 | n32750_o;
  /* divider.vhdl:81:33  */
  assign n32752_o = dend[127:0];
  /* divider.vhdl:81:48  */
  assign n32754_o = {n32752_o, 1'b0};
  /* divider.vhdl:82:33  */
  assign n32755_o = quot[62:0];
  /* divider.vhdl:82:47  */
  assign n32757_o = {n32755_o, 1'b0};
  /* divider.vhdl:83:36  */
  assign n32759_o = count + 7'b0000001;
  /* divider.vhdl:73:17  */
  assign n32760_o = n32738_o ? n32744_o : n32754_o;
  /* divider.vhdl:73:17  */
  assign n32761_o = n32738_o ? n32747_o : n32757_o;
  /* divider.vhdl:73:17  */
  assign n32762_o = n32738_o ? n32749_o : n32759_o;
  /* divider.vhdl:73:17  */
  assign n32763_o = n32738_o ? n32741_o : n32751_o;
  /* divider.vhdl:67:17  */
  assign n32764_o = n32718_o ? n32726_o : n32760_o;
  /* divider.vhdl:67:17  */
  assign n32765_o = n32718_o ? n32729_o : n32761_o;
  /* divider.vhdl:67:17  */
  assign n32766_o = n32718_o ? n32731_o : n32762_o;
  /* divider.vhdl:67:17  */
  assign n32767_o = n32718_o ? n32720_o : n32763_o;
  /* divider.vhdl:62:13  */
  assign n32768_o = running ? n32764_o : dend;
  /* divider.vhdl:62:13  */
  assign n32769_o = running ? n32765_o : quot;
  /* divider.vhdl:62:13  */
  assign n32770_o = running & n32711_o;
  /* divider.vhdl:62:13  */
  assign n32772_o = running ? n32766_o : 7'b0000000;
  /* divider.vhdl:62:13  */
  assign n32773_o = running ? n32714_o : overflow;
  /* divider.vhdl:62:13  */
  assign n32774_o = running ? n32767_o : ovf32;
  /* divider.vhdl:45:13  */
  assign n32775_o = n32693_o ? n32703_o : n32768_o;
  /* divider.vhdl:45:13  */
  assign n32776_o = n32693_o ? n32704_o : div;
  /* divider.vhdl:45:13  */
  assign n32778_o = n32693_o ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n32769_o;
  /* divider.vhdl:45:13  */
  assign n32780_o = n32693_o ? 1'b1 : n32713_o;
  /* divider.vhdl:45:13  */
  assign n32782_o = n32693_o ? 7'b1111111 : n32772_o;
  /* divider.vhdl:45:13  */
  assign n32783_o = n32693_o ? n32705_o : neg_result;
  /* divider.vhdl:45:13  */
  assign n32784_o = n32693_o ? n32706_o : is_modulus;
  /* divider.vhdl:45:13  */
  assign n32785_o = n32693_o ? n32708_o : is_32bit;
  /* divider.vhdl:45:13  */
  assign n32787_o = n32693_o ? n32709_o : is_signed;
  /* divider.vhdl:45:13  */
  assign n32789_o = n32693_o ? 1'b0 : n32773_o;
  /* divider.vhdl:45:13  */
  assign n32791_o = n32693_o ? 1'b0 : n32774_o;
  /* divider.vhdl:39:13  */
  assign n32793_o = rst ? 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : n32775_o;
  /* divider.vhdl:39:13  */
  assign n32795_o = rst ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n32776_o;
  /* divider.vhdl:39:13  */
  assign n32797_o = rst ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n32778_o;
  /* divider.vhdl:39:13  */
  assign n32799_o = rst ? 1'b0 : n32780_o;
  /* divider.vhdl:39:13  */
  assign n32801_o = rst ? 7'b0000000 : n32782_o;
  /* divider.vhdl:39:13  */
  assign n32802_o = rst ? neg_result : n32783_o;
  /* divider.vhdl:39:13  */
  assign n32803_o = rst ? is_modulus : n32784_o;
  /* divider.vhdl:39:13  */
  assign n32804_o = rst ? is_32bit : n32785_o;
  /* divider.vhdl:39:13  */
  assign n32806_o = rst ? is_signed : n32787_o;
  /* divider.vhdl:39:13  */
  assign n32807_o = rst ? overflow : n32789_o;
  /* divider.vhdl:39:13  */
  assign n32808_o = rst ? ovf32 : n32791_o;
  /* divider.vhdl:94:27  */
  assign n32823_o = dend[128:65];
  /* divider.vhdl:93:9  */
  assign n32824_o = is_modulus ? n32823_o : quot;
  /* divider.vhdl:99:55  */
  assign n32826_o = {1'b0, result};
  /* divider.vhdl:99:42  */
  assign n32827_o = -n32826_o;
  /* divider.vhdl:101:28  */
  assign n32829_o = {1'b0, result};
  /* divider.vhdl:98:9  */
  assign n32830_o = neg_result ? n32827_o : n32829_o;
  /* divider.vhdl:104:21  */
  assign n32831_o = ~is_32bit;
  /* divider.vhdl:105:59  */
  assign n32832_o = sresult[64];
  /* divider.vhdl:105:75  */
  assign n32833_o = sresult[63];
  /* divider.vhdl:105:64  */
  assign n32834_o = n32832_o ^ n32833_o;
  /* divider.vhdl:105:47  */
  assign n32835_o = is_signed & n32834_o;
  /* divider.vhdl:105:33  */
  assign n32836_o = overflow | n32835_o;
  /* divider.vhdl:107:38  */
  assign n32837_o = sresult[32];
  /* divider.vhdl:107:53  */
  assign n32838_o = sresult[31];
  /* divider.vhdl:107:43  */
  assign n32839_o = n32837_o != n32838_o;
  /* divider.vhdl:107:28  */
  assign n32840_o = ovf32 | n32839_o;
  /* divider.vhdl:107:13  */
  assign n32843_o = n32840_o ? 1'b1 : 1'b0;
  /* divider.vhdl:106:9  */
  assign n32844_o = is_signed ? n32843_o : ovf32;
  /* divider.vhdl:104:9  */
  assign n32845_o = n32831_o ? n32836_o : n32844_o;
  /* divider.vhdl:115:48  */
  assign n32847_o = ~is_modulus;
  /* divider.vhdl:115:32  */
  assign n32848_o = is_32bit & n32847_o;
  /* divider.vhdl:117:45  */
  assign n32849_o = sresult[31:0];
  /* divider.vhdl:117:36  */
  assign n32851_o = {32'b00000000000000000000000000000000, n32849_o};
  /* divider.vhdl:119:31  */
  assign n32852_o = sresult[63:0];
  /* divider.vhdl:115:9  */
  assign n32853_o = n32848_o ? n32851_o : n32852_o;
  /* divider.vhdl:113:9  */
  assign n32855_o = did_ovf ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n32853_o;
  /* divider.vhdl:129:22  */
  assign n32861_o = count == 7'b1000000;
  /* divider.vhdl:129:13  */
  assign n32863_o = n32861_o ? 1'b1 : 1'b0;
  assign n32864_o = {did_ovf, oresult, n32863_o};
  /* divider.vhdl:38:9  */
  always @(posedge clk)
    n32867_q <= n32793_o;
  /* divider.vhdl:38:9  */
  always @(posedge clk)
    n32868_q <= n32795_o;
  /* divider.vhdl:38:9  */
  always @(posedge clk)
    n32869_q <= n32797_o;
  /* divider.vhdl:38:9  */
  always @(posedge clk)
    n32870_q <= n32799_o;
  /* divider.vhdl:38:9  */
  always @(posedge clk)
    n32871_q <= n32801_o;
  /* divider.vhdl:38:9  */
  always @(posedge clk)
    n32872_q <= n32802_o;
  /* divider.vhdl:38:9  */
  always @(posedge clk)
    n32873_q <= n32803_o;
  /* divider.vhdl:38:9  */
  always @(posedge clk)
    n32874_q <= n32804_o;
  /* divider.vhdl:38:9  */
  always @(posedge clk)
    n32876_q <= n32806_o;
  /* divider.vhdl:38:9  */
  always @(posedge clk)
    n32877_q <= n32807_o;
  /* divider.vhdl:38:9  */
  always @(posedge clk)
    n32878_q <= n32808_o;
  /* divider.vhdl:125:9  */
  always @(posedge clk)
    n32879_q <= n32864_o;
endmodule

module multiply_2
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  clk,
   input  m_in_valid,
   input  [63:0] m_in_data1,
   input  [63:0] m_in_data2,
   input  [127:0] m_in_addend,
   input  m_in_is_32bit,
   input  m_in_not_result,
   output m_out_valid,
   output [127:0] m_out_result,
   output m_out_overflow);
  wire [258:0] n32622_o;
  wire n32624_o;
  wire [127:0] n32625_o;
  wire n32626_o;
  reg [258:0] m;
  reg [5:0] r;
  reg [5:0] rin;
  wire overflow;
  wire ovf_in;
  wire [127:0] mult_out;
  wire [127:0] multiplier_o;
  wire [63:0] n32636_o;
  wire [63:0] n32637_o;
  wire [127:0] n32638_o;
  wire n32645_o;
  wire n32648_o;
  wire n32650_o;
  wire [2:0] n32651_o;
  wire [5:0] n32652_o;
  wire [2:0] n32653_o;
  wire n32654_o;
  wire [127:0] n32655_o;
  wire [127:0] n32656_o;
  wire [5:0] n32657_o;
  wire [2:0] n32658_o;
  wire n32659_o;
  wire [32:0] n32660_o;
  wire n32661_o;
  wire [32:0] n32662_o;
  wire n32663_o;
  wire n32664_o;
  wire n32665_o;
  wire [64:0] n32666_o;
  wire n32667_o;
  wire [64:0] n32668_o;
  wire n32669_o;
  wire n32670_o;
  wire n32671_o;
  wire n32672_o;
  wire [5:0] n32674_o;
  wire [2:0] n32675_o;
  wire n32676_o;
  wire [5:0] n32677_o;
  reg [258:0] n32682_q;
  reg [5:0] n32683_q;
  reg n32684_q;
  wire [129:0] n32685_o;
  assign m_out_valid = n32624_o;
  assign m_out_result = n32625_o;
  assign m_out_overflow = n32626_o;
  assign n32622_o = {m_in_not_result, m_in_is_32bit, m_in_addend, m_in_data2, m_in_data1, m_in_valid};
  assign n32624_o = n32685_o[0];
  assign n32625_o = n32685_o[128:1];
  assign n32626_o = n32685_o[129];
  /* asic/multiply.vhdl:21:12  */
  always @*
    m = n32682_q; // (isignal)
  initial
    m = 259'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* asic/multiply.vhdl:39:12  */
  always @*
    r = n32683_q; // (isignal)
  initial
    r = 6'b000000;
  /* asic/multiply.vhdl:39:15  */
  always @*
    rin = n32677_o; // (isignal)
  initial
    rin = 6'b000000;
  /* asic/multiply.vhdl:40:12  */
  assign overflow = n32684_q; // (signal)
  /* asic/multiply.vhdl:41:12  */
  assign ovf_in = n32672_o; // (signal)
  /* asic/multiply.vhdl:43:12  */
  assign mult_out = multiplier_o; // (signal)
  /* asic/multiply.vhdl:63:5  */
  multiply_add_64x64 multiplier (
`ifdef USE_POWER_PINS
    .VPWR(vccd1),
    .VGND(vssd1),
`endif
    .clk(clk),
    .a(n32636_o),
    .b(n32637_o),
    .c(n32638_o),
    .o(multiplier_o));
  /* asic/multiply.vhdl:66:20  */
  assign n32636_o = m[64:1];
  /* asic/multiply.vhdl:67:20  */
  assign n32637_o = m[128:65];
  /* asic/multiply.vhdl:68:20  */
  assign n32638_o = m[256:129];
  /* asic/multiply.vhdl:79:43  */
  assign n32645_o = m[0];
  /* asic/multiply.vhdl:80:46  */
  assign n32648_o = m[257];
  /* asic/multiply.vhdl:81:45  */
  assign n32650_o = m[258];
  /* asic/multiply.vhdl:84:58  */
  assign n32651_o = r[5:3];
  assign n32652_o = {n32650_o, n32648_o, n32645_o, n32651_o};
  /* asic/multiply.vhdl:87:31  */
  assign n32653_o = n32652_o[2:0];
  /* asic/multiply.vhdl:87:50  */
  assign n32654_o = n32653_o[2];
  /* asic/multiply.vhdl:88:18  */
  assign n32655_o = ~mult_out;
  /* asic/multiply.vhdl:87:9  */
  assign n32656_o = n32654_o ? n32655_o : mult_out;
  assign n32657_o = {n32650_o, n32648_o, n32645_o, n32651_o};
  /* asic/multiply.vhdl:94:31  */
  assign n32658_o = n32657_o[2:0];
  /* asic/multiply.vhdl:94:50  */
  assign n32659_o = n32658_o[1];
  /* asic/multiply.vhdl:95:24  */
  assign n32660_o = n32656_o[63:31];
  /* asic/multiply.vhdl:95:20  */
  assign n32661_o = |(n32660_o);
  /* asic/multiply.vhdl:95:54  */
  assign n32662_o = n32656_o[63:31];
  /* asic/multiply.vhdl:95:49  */
  assign n32663_o = &(n32662_o);
  /* asic/multiply.vhdl:95:44  */
  assign n32664_o = ~n32663_o;
  /* asic/multiply.vhdl:95:40  */
  assign n32665_o = n32661_o & n32664_o;
  /* asic/multiply.vhdl:97:24  */
  assign n32666_o = n32656_o[127:63];
  /* asic/multiply.vhdl:97:20  */
  assign n32667_o = |(n32666_o);
  /* asic/multiply.vhdl:97:55  */
  assign n32668_o = n32656_o[127:63];
  /* asic/multiply.vhdl:97:50  */
  assign n32669_o = &(n32668_o);
  /* asic/multiply.vhdl:97:45  */
  assign n32670_o = ~n32669_o;
  /* asic/multiply.vhdl:97:41  */
  assign n32671_o = n32667_o & n32670_o;
  /* asic/multiply.vhdl:94:9  */
  assign n32672_o = n32659_o ? n32665_o : n32671_o;
  assign n32674_o = {n32650_o, n32648_o, n32645_o, n32651_o};
  /* asic/multiply.vhdl:103:43  */
  assign n32675_o = n32674_o[2:0];
  /* asic/multiply.vhdl:103:62  */
  assign n32676_o = n32675_o[0];
  assign n32677_o = {n32650_o, n32648_o, n32645_o, n32651_o};
  /* asic/multiply.vhdl:56:9  */
  always @(posedge clk)
    n32682_q <= n32622_o;
  initial
    n32682_q = 259'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* asic/multiply.vhdl:56:9  */
  always @(posedge clk)
    n32683_q <= rin;
  initial
    n32683_q = 6'b000000;
  /* asic/multiply.vhdl:56:9  */
  always @(posedge clk)
    n32684_q <= ovf_in;
  /* asic/multiply.vhdl:56:9  */
  assign n32685_o = {overflow, n32656_o, n32676_o};
endmodule

module bit_counter
  (input  clk,
   input  [63:0] rs,
   input  count_right,
   input  do_popcnt,
   input  is_32bit,
   input  [3:0] datalen,
   output [63:0] result);
  wire [63:0] inp;
  wire [63:0] inp_r;
  wire [64:0] sum;
  wire [64:0] sum_r;
  wire [63:0] onehot;
  wire [63:0] \edge ;
  wire [5:0] bitnum;
  wire [63:0] cntz;
  wire [3:0] dlen_r;
  wire pcnt_r;
  wire [63:0] pc2;
  wire [47:0] pc4;
  wire [31:0] pc8;
  wire [31:0] pc8_r;
  wire [11:0] pc32;
  wire [63:0] popcnt;
  wire n31308_o;
  wire n31309_o;
  wire n31316_o;
  wire n31319_o;
  wire n31321_o;
  wire n31323_o;
  wire n31325_o;
  wire n31327_o;
  wire n31329_o;
  wire n31331_o;
  wire n31333_o;
  wire n31335_o;
  wire n31337_o;
  wire n31339_o;
  wire n31341_o;
  wire n31343_o;
  wire n31345_o;
  wire n31347_o;
  wire n31349_o;
  wire n31351_o;
  wire n31353_o;
  wire n31355_o;
  wire n31357_o;
  wire n31359_o;
  wire n31361_o;
  wire n31363_o;
  wire n31365_o;
  wire n31367_o;
  wire n31369_o;
  wire n31371_o;
  wire n31373_o;
  wire n31375_o;
  wire n31377_o;
  wire n31379_o;
  wire n31381_o;
  wire n31383_o;
  wire n31385_o;
  wire n31387_o;
  wire n31389_o;
  wire n31391_o;
  wire n31393_o;
  wire n31395_o;
  wire n31397_o;
  wire n31399_o;
  wire n31401_o;
  wire n31403_o;
  wire n31405_o;
  wire n31407_o;
  wire n31409_o;
  wire n31411_o;
  wire n31413_o;
  wire n31415_o;
  wire n31417_o;
  wire n31419_o;
  wire n31421_o;
  wire n31423_o;
  wire n31425_o;
  wire n31427_o;
  wire n31429_o;
  wire n31431_o;
  wire n31433_o;
  wire n31435_o;
  wire n31437_o;
  wire n31439_o;
  wire n31441_o;
  wire n31443_o;
  wire [63:0] n31444_o;
  wire [63:0] n31445_o;
  wire n31447_o;
  wire [31:0] n31449_o;
  wire n31455_o;
  wire n31458_o;
  wire n31460_o;
  wire n31462_o;
  wire n31464_o;
  wire n31466_o;
  wire n31468_o;
  wire n31470_o;
  wire n31472_o;
  wire n31474_o;
  wire n31476_o;
  wire n31478_o;
  wire n31480_o;
  wire n31482_o;
  wire n31484_o;
  wire n31486_o;
  wire n31488_o;
  wire n31490_o;
  wire n31492_o;
  wire n31494_o;
  wire n31496_o;
  wire n31498_o;
  wire n31500_o;
  wire n31502_o;
  wire n31504_o;
  wire n31506_o;
  wire n31508_o;
  wire n31510_o;
  wire n31512_o;
  wire n31514_o;
  wire n31516_o;
  wire n31518_o;
  wire [31:0] n31519_o;
  wire [31:0] n31520_o;
  wire [31:0] n31521_o;
  wire [63:0] n31522_o;
  wire [63:0] n31523_o;
  wire [63:0] n31524_o;
  wire [64:0] n31526_o;
  wire [64:0] n31528_o;
  wire [63:0] n31529_o;
  wire [63:0] n31530_o;
  wire n31540_o;
  wire n31541_o;
  wire n31542_o;
  wire n31543_o;
  wire n31545_o;
  wire n31547_o;
  wire n31548_o;
  wire n31549_o;
  wire n31550_o;
  wire n31551_o;
  wire n31552_o;
  wire n31553_o;
  wire n31554_o;
  wire n31555_o;
  wire n31556_o;
  wire n31557_o;
  wire n31558_o;
  wire n31559_o;
  wire n31560_o;
  wire n31561_o;
  wire n31562_o;
  wire n31563_o;
  wire n31564_o;
  wire n31565_o;
  wire n31566_o;
  wire n31567_o;
  wire n31568_o;
  wire n31569_o;
  wire n31570_o;
  wire n31571_o;
  wire n31572_o;
  wire n31573_o;
  wire n31574_o;
  wire n31575_o;
  wire n31576_o;
  wire n31577_o;
  wire n31578_o;
  wire n31579_o;
  wire n31580_o;
  wire n31581_o;
  wire n31582_o;
  wire n31583_o;
  wire n31584_o;
  wire n31585_o;
  wire n31586_o;
  wire n31587_o;
  wire n31588_o;
  wire n31589_o;
  wire n31590_o;
  wire n31591_o;
  wire n31592_o;
  wire n31593_o;
  wire n31594_o;
  wire n31595_o;
  wire n31596_o;
  wire n31597_o;
  wire n31598_o;
  wire n31599_o;
  wire n31600_o;
  wire n31601_o;
  wire n31602_o;
  wire n31603_o;
  wire n31604_o;
  wire n31605_o;
  wire n31606_o;
  wire n31607_o;
  wire n31608_o;
  wire n31609_o;
  wire n31610_o;
  wire n31611_o;
  wire n31612_o;
  wire n31613_o;
  wire n31614_o;
  wire n31615_o;
  wire n31616_o;
  wire n31617_o;
  wire n31618_o;
  wire n31619_o;
  wire n31620_o;
  wire n31621_o;
  wire n31622_o;
  wire n31623_o;
  wire n31624_o;
  wire n31625_o;
  wire n31626_o;
  wire n31627_o;
  wire n31628_o;
  wire n31629_o;
  wire n31630_o;
  wire n31631_o;
  wire n31632_o;
  wire n31633_o;
  wire n31634_o;
  wire n31635_o;
  wire n31636_o;
  wire n31637_o;
  wire n31638_o;
  wire n31639_o;
  wire n31640_o;
  wire n31641_o;
  wire n31642_o;
  wire n31643_o;
  wire n31644_o;
  wire n31645_o;
  wire n31646_o;
  wire n31647_o;
  wire n31648_o;
  wire n31649_o;
  wire n31650_o;
  wire n31651_o;
  wire n31652_o;
  wire n31653_o;
  wire n31654_o;
  wire n31655_o;
  wire n31656_o;
  wire n31657_o;
  wire n31658_o;
  wire n31659_o;
  wire n31660_o;
  wire n31661_o;
  wire n31662_o;
  wire n31663_o;
  wire n31664_o;
  wire n31665_o;
  wire n31666_o;
  wire n31667_o;
  wire n31668_o;
  wire n31669_o;
  wire n31670_o;
  wire n31671_o;
  wire n31672_o;
  wire n31673_o;
  wire n31674_o;
  wire n31675_o;
  wire n31676_o;
  wire n31677_o;
  wire n31678_o;
  wire n31679_o;
  wire n31680_o;
  wire n31681_o;
  wire n31682_o;
  wire n31683_o;
  wire n31684_o;
  wire n31685_o;
  wire n31686_o;
  wire n31687_o;
  wire n31688_o;
  wire n31689_o;
  wire n31690_o;
  wire n31691_o;
  wire n31692_o;
  wire n31693_o;
  wire n31694_o;
  wire n31695_o;
  wire n31696_o;
  wire n31697_o;
  wire n31698_o;
  wire n31699_o;
  wire n31700_o;
  wire n31701_o;
  wire n31704_o;
  wire n31705_o;
  wire n31706_o;
  wire n31707_o;
  wire n31709_o;
  wire n31711_o;
  wire n31712_o;
  wire n31713_o;
  wire n31714_o;
  wire n31715_o;
  wire n31716_o;
  wire n31717_o;
  wire n31718_o;
  wire n31719_o;
  wire n31720_o;
  wire n31721_o;
  wire n31722_o;
  wire n31723_o;
  wire n31724_o;
  wire n31725_o;
  wire n31726_o;
  wire n31727_o;
  wire n31728_o;
  wire n31729_o;
  wire n31730_o;
  wire n31731_o;
  wire n31732_o;
  wire n31733_o;
  wire n31734_o;
  wire n31735_o;
  wire n31736_o;
  wire n31737_o;
  wire n31738_o;
  wire n31739_o;
  wire n31740_o;
  wire n31741_o;
  wire n31742_o;
  wire n31743_o;
  wire n31744_o;
  wire n31745_o;
  wire n31746_o;
  wire n31747_o;
  wire n31748_o;
  wire n31749_o;
  wire n31750_o;
  wire n31751_o;
  wire n31752_o;
  wire n31753_o;
  wire n31754_o;
  wire n31755_o;
  wire n31756_o;
  wire n31757_o;
  wire n31758_o;
  wire n31759_o;
  wire n31760_o;
  wire n31761_o;
  wire n31762_o;
  wire n31763_o;
  wire n31764_o;
  wire n31765_o;
  wire n31766_o;
  wire n31767_o;
  wire n31768_o;
  wire n31769_o;
  wire n31770_o;
  wire n31771_o;
  wire n31772_o;
  wire n31773_o;
  wire n31774_o;
  wire n31775_o;
  wire n31776_o;
  wire n31777_o;
  wire n31778_o;
  wire n31779_o;
  wire n31780_o;
  wire n31781_o;
  wire n31782_o;
  wire n31783_o;
  wire n31784_o;
  wire n31785_o;
  wire n31787_o;
  wire n31788_o;
  wire n31789_o;
  wire n31790_o;
  wire n31792_o;
  wire n31794_o;
  wire n31795_o;
  wire n31796_o;
  wire n31797_o;
  wire n31798_o;
  wire n31799_o;
  wire n31800_o;
  wire n31801_o;
  wire n31802_o;
  wire n31803_o;
  wire n31804_o;
  wire n31805_o;
  wire n31806_o;
  wire n31807_o;
  wire n31808_o;
  wire n31809_o;
  wire n31810_o;
  wire n31811_o;
  wire n31812_o;
  wire n31813_o;
  wire n31814_o;
  wire n31815_o;
  wire n31816_o;
  wire n31817_o;
  wire n31818_o;
  wire n31819_o;
  wire n31820_o;
  wire n31821_o;
  wire n31822_o;
  wire n31823_o;
  wire n31824_o;
  wire n31825_o;
  wire n31826_o;
  wire n31827_o;
  wire n31828_o;
  wire n31830_o;
  wire n31831_o;
  wire n31832_o;
  wire n31833_o;
  wire n31835_o;
  wire n31837_o;
  wire n31838_o;
  wire n31839_o;
  wire n31840_o;
  wire n31841_o;
  wire n31842_o;
  wire n31843_o;
  wire n31844_o;
  wire n31845_o;
  wire n31846_o;
  wire n31847_o;
  wire n31848_o;
  wire n31849_o;
  wire n31850_o;
  wire n31851_o;
  wire n31853_o;
  wire n31854_o;
  wire n31855_o;
  wire n31856_o;
  wire n31858_o;
  wire n31860_o;
  wire n31861_o;
  wire n31862_o;
  wire n31863_o;
  wire n31864_o;
  wire n31866_o;
  wire n31867_o;
  wire n31868_o;
  wire n31869_o;
  wire n31871_o;
  wire [5:0] n31873_o;
  wire [63:0] n31874_o;
  wire [63:0] n31875_o;
  wire n31885_o;
  wire n31886_o;
  wire n31888_o;
  wire n31890_o;
  wire n31891_o;
  wire n31892_o;
  wire n31893_o;
  wire n31894_o;
  wire n31895_o;
  wire n31896_o;
  wire n31897_o;
  wire n31898_o;
  wire n31899_o;
  wire n31900_o;
  wire n31901_o;
  wire n31902_o;
  wire n31903_o;
  wire n31904_o;
  wire n31905_o;
  wire n31906_o;
  wire n31907_o;
  wire n31908_o;
  wire n31909_o;
  wire n31910_o;
  wire n31911_o;
  wire n31912_o;
  wire n31913_o;
  wire n31914_o;
  wire n31915_o;
  wire n31916_o;
  wire n31917_o;
  wire n31918_o;
  wire n31919_o;
  wire n31920_o;
  wire n31921_o;
  wire n31922_o;
  wire n31923_o;
  wire n31924_o;
  wire n31925_o;
  wire n31926_o;
  wire n31927_o;
  wire n31928_o;
  wire n31929_o;
  wire n31930_o;
  wire n31931_o;
  wire n31932_o;
  wire n31933_o;
  wire n31934_o;
  wire n31935_o;
  wire n31936_o;
  wire n31937_o;
  wire n31938_o;
  wire n31939_o;
  wire n31940_o;
  wire n31941_o;
  wire n31942_o;
  wire n31943_o;
  wire n31944_o;
  wire n31945_o;
  wire n31946_o;
  wire n31947_o;
  wire n31948_o;
  wire n31949_o;
  wire n31950_o;
  wire n31951_o;
  wire n31952_o;
  wire n31953_o;
  wire n31954_o;
  wire n31955_o;
  wire n31956_o;
  wire n31957_o;
  wire n31958_o;
  wire n31959_o;
  wire n31960_o;
  wire n31961_o;
  wire n31962_o;
  wire n31963_o;
  wire n31964_o;
  wire n31965_o;
  wire n31966_o;
  wire n31967_o;
  wire n31968_o;
  wire n31969_o;
  wire n31970_o;
  wire n31971_o;
  wire n31972_o;
  wire n31973_o;
  wire n31974_o;
  wire n31975_o;
  wire n31976_o;
  wire n31977_o;
  wire n31978_o;
  wire n31979_o;
  wire n31980_o;
  wire n31981_o;
  wire n31982_o;
  wire [1:0] n31985_o;
  wire n31986_o;
  wire n31988_o;
  wire [1:0] n31990_o;
  wire n31991_o;
  wire n31992_o;
  wire [1:0] n31993_o;
  wire n31994_o;
  wire n31995_o;
  wire [1:0] n31996_o;
  wire n31997_o;
  wire n31998_o;
  wire [1:0] n31999_o;
  wire n32000_o;
  wire n32001_o;
  wire [1:0] n32002_o;
  wire n32003_o;
  wire n32004_o;
  wire [1:0] n32005_o;
  wire n32006_o;
  wire n32007_o;
  wire [1:0] n32008_o;
  wire n32009_o;
  wire n32010_o;
  wire [1:0] n32011_o;
  wire n32012_o;
  wire n32013_o;
  wire [1:0] n32014_o;
  wire n32015_o;
  wire n32016_o;
  wire [1:0] n32017_o;
  wire n32018_o;
  wire n32019_o;
  wire [1:0] n32020_o;
  wire n32021_o;
  wire n32022_o;
  wire [1:0] n32023_o;
  wire n32024_o;
  wire n32025_o;
  wire [1:0] n32026_o;
  wire n32027_o;
  wire n32028_o;
  wire [1:0] n32029_o;
  wire n32030_o;
  wire n32031_o;
  wire [1:0] n32032_o;
  wire n32033_o;
  wire n32034_o;
  wire [3:0] n32036_o;
  wire n32037_o;
  wire n32039_o;
  wire [3:0] n32041_o;
  wire n32042_o;
  wire n32043_o;
  wire [3:0] n32044_o;
  wire n32045_o;
  wire n32046_o;
  wire [3:0] n32047_o;
  wire n32048_o;
  wire n32049_o;
  wire [3:0] n32050_o;
  wire n32051_o;
  wire n32052_o;
  wire [3:0] n32053_o;
  wire n32054_o;
  wire n32055_o;
  wire [3:0] n32056_o;
  wire n32057_o;
  wire n32058_o;
  wire [3:0] n32059_o;
  wire n32060_o;
  wire n32061_o;
  wire [7:0] n32063_o;
  wire n32064_o;
  wire n32066_o;
  wire [7:0] n32068_o;
  wire n32069_o;
  wire n32070_o;
  wire [7:0] n32071_o;
  wire n32072_o;
  wire n32073_o;
  wire [7:0] n32074_o;
  wire n32075_o;
  wire n32076_o;
  wire [15:0] n32078_o;
  wire n32079_o;
  wire n32081_o;
  wire [15:0] n32083_o;
  wire n32084_o;
  wire n32085_o;
  wire [31:0] n32087_o;
  wire n32088_o;
  wire n32090_o;
  wire [5:0] n32092_o;
  wire [3:0] n32093_o;
  wire [1:0] n32094_o;
  wire n32095_o;
  wire [57:0] n32097_o;
  wire [63:0] n32098_o;
  wire [3:0] n32102_o;
  wire [3:0] n32103_o;
  wire [3:0] n32104_o;
  wire [3:0] n32105_o;
  wire [3:0] n32106_o;
  wire [3:0] n32107_o;
  wire [3:0] n32108_o;
  wire [3:0] n32109_o;
  wire [31:0] n32112_o;
  wire n32116_o;
  wire [1:0] n32118_o;
  wire n32119_o;
  wire [1:0] n32121_o;
  wire [1:0] n32122_o;
  wire n32123_o;
  wire [1:0] n32125_o;
  wire n32126_o;
  wire [1:0] n32128_o;
  wire [1:0] n32129_o;
  wire n32130_o;
  wire [1:0] n32132_o;
  wire n32133_o;
  wire [1:0] n32135_o;
  wire [1:0] n32136_o;
  wire n32137_o;
  wire [1:0] n32139_o;
  wire n32140_o;
  wire [1:0] n32142_o;
  wire [1:0] n32143_o;
  wire n32144_o;
  wire [1:0] n32146_o;
  wire n32147_o;
  wire [1:0] n32149_o;
  wire [1:0] n32150_o;
  wire n32151_o;
  wire [1:0] n32153_o;
  wire n32154_o;
  wire [1:0] n32156_o;
  wire [1:0] n32157_o;
  wire n32158_o;
  wire [1:0] n32160_o;
  wire n32161_o;
  wire [1:0] n32163_o;
  wire [1:0] n32164_o;
  wire n32165_o;
  wire [1:0] n32167_o;
  wire n32168_o;
  wire [1:0] n32170_o;
  wire [1:0] n32171_o;
  wire n32172_o;
  wire [1:0] n32174_o;
  wire n32175_o;
  wire [1:0] n32177_o;
  wire [1:0] n32178_o;
  wire n32179_o;
  wire [1:0] n32181_o;
  wire n32182_o;
  wire [1:0] n32184_o;
  wire [1:0] n32185_o;
  wire n32186_o;
  wire [1:0] n32188_o;
  wire n32189_o;
  wire [1:0] n32191_o;
  wire [1:0] n32192_o;
  wire n32193_o;
  wire [1:0] n32195_o;
  wire n32196_o;
  wire [1:0] n32198_o;
  wire [1:0] n32199_o;
  wire n32200_o;
  wire [1:0] n32202_o;
  wire n32203_o;
  wire [1:0] n32205_o;
  wire [1:0] n32206_o;
  wire n32207_o;
  wire [1:0] n32209_o;
  wire n32210_o;
  wire [1:0] n32212_o;
  wire [1:0] n32213_o;
  wire n32214_o;
  wire [1:0] n32216_o;
  wire n32217_o;
  wire [1:0] n32219_o;
  wire [1:0] n32220_o;
  wire n32221_o;
  wire [1:0] n32223_o;
  wire n32224_o;
  wire [1:0] n32226_o;
  wire [1:0] n32227_o;
  wire n32228_o;
  wire [1:0] n32230_o;
  wire n32231_o;
  wire [1:0] n32233_o;
  wire [1:0] n32234_o;
  wire n32235_o;
  wire [1:0] n32237_o;
  wire n32238_o;
  wire [1:0] n32240_o;
  wire [1:0] n32241_o;
  wire n32242_o;
  wire [1:0] n32244_o;
  wire n32245_o;
  wire [1:0] n32247_o;
  wire [1:0] n32248_o;
  wire n32249_o;
  wire [1:0] n32251_o;
  wire n32252_o;
  wire [1:0] n32254_o;
  wire [1:0] n32255_o;
  wire n32256_o;
  wire [1:0] n32258_o;
  wire n32259_o;
  wire [1:0] n32261_o;
  wire [1:0] n32262_o;
  wire n32263_o;
  wire [1:0] n32265_o;
  wire n32266_o;
  wire [1:0] n32268_o;
  wire [1:0] n32269_o;
  wire n32270_o;
  wire [1:0] n32272_o;
  wire n32273_o;
  wire [1:0] n32275_o;
  wire [1:0] n32276_o;
  wire n32277_o;
  wire [1:0] n32279_o;
  wire n32280_o;
  wire [1:0] n32282_o;
  wire [1:0] n32283_o;
  wire n32284_o;
  wire [1:0] n32286_o;
  wire n32287_o;
  wire [1:0] n32289_o;
  wire [1:0] n32290_o;
  wire n32291_o;
  wire [1:0] n32293_o;
  wire n32294_o;
  wire [1:0] n32296_o;
  wire [1:0] n32297_o;
  wire n32298_o;
  wire [1:0] n32300_o;
  wire n32301_o;
  wire [1:0] n32303_o;
  wire [1:0] n32304_o;
  wire n32305_o;
  wire [1:0] n32307_o;
  wire n32308_o;
  wire [1:0] n32310_o;
  wire [1:0] n32311_o;
  wire n32312_o;
  wire [1:0] n32314_o;
  wire n32315_o;
  wire [1:0] n32317_o;
  wire [1:0] n32318_o;
  wire n32319_o;
  wire [1:0] n32321_o;
  wire n32322_o;
  wire [1:0] n32324_o;
  wire [1:0] n32325_o;
  wire n32326_o;
  wire [1:0] n32328_o;
  wire n32329_o;
  wire [1:0] n32331_o;
  wire [1:0] n32332_o;
  wire n32333_o;
  wire [1:0] n32335_o;
  wire n32336_o;
  wire [1:0] n32338_o;
  wire [1:0] n32339_o;
  wire [1:0] n32340_o;
  wire [2:0] n32342_o;
  wire [1:0] n32343_o;
  wire [2:0] n32345_o;
  wire [2:0] n32346_o;
  wire [1:0] n32347_o;
  wire [2:0] n32349_o;
  wire [1:0] n32350_o;
  wire [2:0] n32352_o;
  wire [2:0] n32353_o;
  wire [1:0] n32354_o;
  wire [2:0] n32356_o;
  wire [1:0] n32357_o;
  wire [2:0] n32359_o;
  wire [2:0] n32360_o;
  wire [1:0] n32361_o;
  wire [2:0] n32363_o;
  wire [1:0] n32364_o;
  wire [2:0] n32366_o;
  wire [2:0] n32367_o;
  wire [1:0] n32368_o;
  wire [2:0] n32370_o;
  wire [1:0] n32371_o;
  wire [2:0] n32373_o;
  wire [2:0] n32374_o;
  wire [1:0] n32375_o;
  wire [2:0] n32377_o;
  wire [1:0] n32378_o;
  wire [2:0] n32380_o;
  wire [2:0] n32381_o;
  wire [1:0] n32382_o;
  wire [2:0] n32384_o;
  wire [1:0] n32385_o;
  wire [2:0] n32387_o;
  wire [2:0] n32388_o;
  wire [1:0] n32389_o;
  wire [2:0] n32391_o;
  wire [1:0] n32392_o;
  wire [2:0] n32394_o;
  wire [2:0] n32395_o;
  wire [1:0] n32396_o;
  wire [2:0] n32398_o;
  wire [1:0] n32399_o;
  wire [2:0] n32401_o;
  wire [2:0] n32402_o;
  wire [1:0] n32403_o;
  wire [2:0] n32405_o;
  wire [1:0] n32406_o;
  wire [2:0] n32408_o;
  wire [2:0] n32409_o;
  wire [1:0] n32410_o;
  wire [2:0] n32412_o;
  wire [1:0] n32413_o;
  wire [2:0] n32415_o;
  wire [2:0] n32416_o;
  wire [1:0] n32417_o;
  wire [2:0] n32419_o;
  wire [1:0] n32420_o;
  wire [2:0] n32422_o;
  wire [2:0] n32423_o;
  wire [1:0] n32424_o;
  wire [2:0] n32426_o;
  wire [1:0] n32427_o;
  wire [2:0] n32429_o;
  wire [2:0] n32430_o;
  wire [1:0] n32431_o;
  wire [2:0] n32433_o;
  wire [1:0] n32434_o;
  wire [2:0] n32436_o;
  wire [2:0] n32437_o;
  wire [1:0] n32438_o;
  wire [2:0] n32440_o;
  wire [1:0] n32441_o;
  wire [2:0] n32443_o;
  wire [2:0] n32444_o;
  wire [1:0] n32445_o;
  wire [2:0] n32447_o;
  wire [1:0] n32448_o;
  wire [2:0] n32450_o;
  wire [2:0] n32451_o;
  wire [2:0] n32452_o;
  wire [3:0] n32454_o;
  wire [2:0] n32455_o;
  wire [3:0] n32457_o;
  wire [3:0] n32458_o;
  wire [2:0] n32459_o;
  wire [3:0] n32461_o;
  wire [2:0] n32462_o;
  wire [3:0] n32464_o;
  wire [3:0] n32465_o;
  wire [2:0] n32466_o;
  wire [3:0] n32468_o;
  wire [2:0] n32469_o;
  wire [3:0] n32471_o;
  wire [3:0] n32472_o;
  wire [2:0] n32473_o;
  wire [3:0] n32475_o;
  wire [2:0] n32476_o;
  wire [3:0] n32478_o;
  wire [3:0] n32479_o;
  wire [2:0] n32480_o;
  wire [3:0] n32482_o;
  wire [2:0] n32483_o;
  wire [3:0] n32485_o;
  wire [3:0] n32486_o;
  wire [2:0] n32487_o;
  wire [3:0] n32489_o;
  wire [2:0] n32490_o;
  wire [3:0] n32492_o;
  wire [3:0] n32493_o;
  wire [2:0] n32494_o;
  wire [3:0] n32496_o;
  wire [2:0] n32497_o;
  wire [3:0] n32499_o;
  wire [3:0] n32500_o;
  wire [2:0] n32501_o;
  wire [3:0] n32503_o;
  wire [2:0] n32504_o;
  wire [3:0] n32506_o;
  wire [3:0] n32507_o;
  wire [3:0] n32508_o;
  wire [5:0] n32510_o;
  wire [3:0] n32511_o;
  wire [5:0] n32513_o;
  wire [5:0] n32514_o;
  wire [3:0] n32515_o;
  wire [5:0] n32517_o;
  wire [5:0] n32518_o;
  wire [3:0] n32519_o;
  wire [5:0] n32521_o;
  wire [5:0] n32522_o;
  wire [3:0] n32523_o;
  wire [5:0] n32525_o;
  wire [3:0] n32526_o;
  wire [5:0] n32528_o;
  wire [5:0] n32529_o;
  wire [3:0] n32530_o;
  wire [5:0] n32532_o;
  wire [5:0] n32533_o;
  wire [3:0] n32534_o;
  wire [5:0] n32536_o;
  wire [5:0] n32537_o;
  wire [1:0] n32538_o;
  wire n32540_o;
  wire [3:0] n32541_o;
  wire [3:0] n32542_o;
  wire [3:0] n32543_o;
  wire [3:0] n32544_o;
  wire [3:0] n32545_o;
  wire [3:0] n32546_o;
  wire [3:0] n32547_o;
  wire [3:0] n32548_o;
  wire n32549_o;
  wire n32550_o;
  wire [5:0] n32551_o;
  wire [5:0] n32552_o;
  wire [5:0] n32553_o;
  wire [6:0] n32555_o;
  wire [5:0] n32556_o;
  wire [6:0] n32558_o;
  wire [6:0] n32559_o;
  wire [5:0] n32560_o;
  wire [5:0] n32561_o;
  wire n32562_o;
  wire n32564_o;
  wire [5:0] n32566_o;
  wire [6:0] n32567_o;
  wire [3:0] n32568_o;
  wire [3:0] n32569_o;
  wire [2:0] n32570_o;
  wire [2:0] n32572_o;
  wire [3:0] n32574_o;
  wire [3:0] n32576_o;
  wire [3:0] n32578_o;
  wire [3:0] n32579_o;
  wire [3:0] n32580_o;
  wire [1:0] n32581_o;
  wire [1:0] n32583_o;
  wire [3:0] n32585_o;
  wire [3:0] n32587_o;
  wire [3:0] n32589_o;
  localparam [63:0] n32590_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire n32594_o;
  wire [3:0] n32596_o;
  wire [3:0] n32598_o;
  wire [3:0] n32600_o;
  wire [1:0] n32603_o;
  wire [3:0] n32605_o;
  wire [3:0] n32606_o;
  wire [3:0] n32607_o;
  wire n32609_o;
  wire [63:0] n32610_o;
  reg [63:0] n32611_q;
  reg [64:0] n32612_q;
  wire [5:0] n32613_o;
  reg [3:0] n32614_q;
  reg n32615_q;
  wire [63:0] n32616_o;
  wire [47:0] n32617_o;
  wire [31:0] n32618_o;
  reg [31:0] n32619_q;
  wire [11:0] n32620_o;
  wire [63:0] n32621_o;
  assign result = n32610_o;
  /* countbits.vhdl:22:12  */
  assign inp = n31523_o; // (signal)
  /* countbits.vhdl:23:12  */
  assign inp_r = n32611_q; // (signal)
  /* countbits.vhdl:24:12  */
  assign sum = n31528_o; // (signal)
  /* countbits.vhdl:25:12  */
  assign sum_r = n32612_q; // (signal)
  /* countbits.vhdl:26:12  */
  assign onehot = n31875_o; // (signal)
  /* countbits.vhdl:27:12  */
  assign \edge  = n31530_o; // (signal)
  /* countbits.vhdl:28:12  */
  assign bitnum = n32613_o; // (signal)
  /* countbits.vhdl:29:12  */
  assign cntz = n32098_o; // (signal)
  /* countbits.vhdl:32:12  */
  assign dlen_r = n32614_q; // (signal)
  /* countbits.vhdl:33:12  */
  assign pcnt_r = n32615_q; // (signal)
  /* countbits.vhdl:36:12  */
  assign pc2 = n32616_o; // (signal)
  /* countbits.vhdl:39:12  */
  assign pc4 = n32617_o; // (signal)
  /* countbits.vhdl:42:12  */
  assign pc8 = n32618_o; // (signal)
  /* countbits.vhdl:43:12  */
  assign pc8_r = n32619_q; // (signal)
  /* countbits.vhdl:46:12  */
  assign pc32 = n32620_o; // (signal)
  /* countbits.vhdl:47:12  */
  assign popcnt = n32621_o; // (signal)
  /* countbits.vhdl:61:21  */
  assign n31308_o = ~is_32bit;
  /* countbits.vhdl:62:28  */
  assign n31309_o = ~count_right;
  /* helpers.vhdl:221:43  */
  assign n31316_o = rs[0];
  /* helpers.vhdl:221:43  */
  assign n31319_o = rs[1];
  /* helpers.vhdl:221:43  */
  assign n31321_o = rs[2];
  /* helpers.vhdl:221:43  */
  assign n31323_o = rs[3];
  /* helpers.vhdl:221:43  */
  assign n31325_o = rs[4];
  /* helpers.vhdl:221:43  */
  assign n31327_o = rs[5];
  /* helpers.vhdl:221:43  */
  assign n31329_o = rs[6];
  /* helpers.vhdl:221:43  */
  assign n31331_o = rs[7];
  /* helpers.vhdl:221:43  */
  assign n31333_o = rs[8];
  /* helpers.vhdl:221:43  */
  assign n31335_o = rs[9];
  /* helpers.vhdl:221:43  */
  assign n31337_o = rs[10];
  /* helpers.vhdl:221:43  */
  assign n31339_o = rs[11];
  /* helpers.vhdl:221:43  */
  assign n31341_o = rs[12];
  /* helpers.vhdl:221:43  */
  assign n31343_o = rs[13];
  /* helpers.vhdl:221:43  */
  assign n31345_o = rs[14];
  /* helpers.vhdl:221:43  */
  assign n31347_o = rs[15];
  /* helpers.vhdl:221:43  */
  assign n31349_o = rs[16];
  /* helpers.vhdl:221:43  */
  assign n31351_o = rs[17];
  /* helpers.vhdl:221:43  */
  assign n31353_o = rs[18];
  /* helpers.vhdl:221:43  */
  assign n31355_o = rs[19];
  /* helpers.vhdl:221:43  */
  assign n31357_o = rs[20];
  /* helpers.vhdl:221:43  */
  assign n31359_o = rs[21];
  /* helpers.vhdl:221:43  */
  assign n31361_o = rs[22];
  /* helpers.vhdl:221:43  */
  assign n31363_o = rs[23];
  /* helpers.vhdl:221:43  */
  assign n31365_o = rs[24];
  /* helpers.vhdl:221:43  */
  assign n31367_o = rs[25];
  /* helpers.vhdl:221:43  */
  assign n31369_o = rs[26];
  /* helpers.vhdl:221:43  */
  assign n31371_o = rs[27];
  /* helpers.vhdl:221:43  */
  assign n31373_o = rs[28];
  /* helpers.vhdl:221:43  */
  assign n31375_o = rs[29];
  /* helpers.vhdl:221:43  */
  assign n31377_o = rs[30];
  /* helpers.vhdl:221:43  */
  assign n31379_o = rs[31];
  /* helpers.vhdl:221:43  */
  assign n31381_o = rs[32];
  /* helpers.vhdl:221:43  */
  assign n31383_o = rs[33];
  /* helpers.vhdl:221:43  */
  assign n31385_o = rs[34];
  /* helpers.vhdl:221:43  */
  assign n31387_o = rs[35];
  /* helpers.vhdl:221:43  */
  assign n31389_o = rs[36];
  /* helpers.vhdl:221:43  */
  assign n31391_o = rs[37];
  /* helpers.vhdl:221:43  */
  assign n31393_o = rs[38];
  /* helpers.vhdl:221:43  */
  assign n31395_o = rs[39];
  /* helpers.vhdl:221:43  */
  assign n31397_o = rs[40];
  /* helpers.vhdl:221:43  */
  assign n31399_o = rs[41];
  /* helpers.vhdl:221:43  */
  assign n31401_o = rs[42];
  /* helpers.vhdl:221:43  */
  assign n31403_o = rs[43];
  /* helpers.vhdl:221:43  */
  assign n31405_o = rs[44];
  /* helpers.vhdl:221:43  */
  assign n31407_o = rs[45];
  /* helpers.vhdl:221:43  */
  assign n31409_o = rs[46];
  /* helpers.vhdl:221:43  */
  assign n31411_o = rs[47];
  /* helpers.vhdl:221:43  */
  assign n31413_o = rs[48];
  /* helpers.vhdl:221:43  */
  assign n31415_o = rs[49];
  /* helpers.vhdl:221:43  */
  assign n31417_o = rs[50];
  /* helpers.vhdl:221:43  */
  assign n31419_o = rs[51];
  /* helpers.vhdl:221:43  */
  assign n31421_o = rs[52];
  /* helpers.vhdl:221:43  */
  assign n31423_o = rs[53];
  /* helpers.vhdl:221:43  */
  assign n31425_o = rs[54];
  /* helpers.vhdl:221:43  */
  assign n31427_o = rs[55];
  /* helpers.vhdl:221:43  */
  assign n31429_o = rs[56];
  /* helpers.vhdl:221:43  */
  assign n31431_o = rs[57];
  /* helpers.vhdl:221:43  */
  assign n31433_o = rs[58];
  /* helpers.vhdl:221:43  */
  assign n31435_o = rs[59];
  /* helpers.vhdl:221:43  */
  assign n31437_o = rs[60];
  /* helpers.vhdl:221:43  */
  assign n31439_o = rs[61];
  /* helpers.vhdl:221:43  */
  assign n31441_o = rs[62];
  /* helpers.vhdl:221:43  */
  assign n31443_o = rs[63];
  assign n31444_o = {n31316_o, n31319_o, n31321_o, n31323_o, n31325_o, n31327_o, n31329_o, n31331_o, n31333_o, n31335_o, n31337_o, n31339_o, n31341_o, n31343_o, n31345_o, n31347_o, n31349_o, n31351_o, n31353_o, n31355_o, n31357_o, n31359_o, n31361_o, n31363_o, n31365_o, n31367_o, n31369_o, n31371_o, n31373_o, n31375_o, n31377_o, n31379_o, n31381_o, n31383_o, n31385_o, n31387_o, n31389_o, n31391_o, n31393_o, n31395_o, n31397_o, n31399_o, n31401_o, n31403_o, n31405_o, n31407_o, n31409_o, n31411_o, n31413_o, n31415_o, n31417_o, n31419_o, n31421_o, n31423_o, n31425_o, n31427_o, n31429_o, n31431_o, n31433_o, n31435_o, n31437_o, n31439_o, n31441_o, n31443_o};
  /* countbits.vhdl:62:13  */
  assign n31445_o = n31309_o ? n31444_o : rs;
  /* countbits.vhdl:69:28  */
  assign n31447_o = ~count_right;
  /* countbits.vhdl:70:51  */
  assign n31449_o = rs[31:0];
  /* helpers.vhdl:221:43  */
  assign n31455_o = n31449_o[0];
  /* helpers.vhdl:221:43  */
  assign n31458_o = n31449_o[1];
  /* helpers.vhdl:221:43  */
  assign n31460_o = n31449_o[2];
  /* helpers.vhdl:221:43  */
  assign n31462_o = n31449_o[3];
  /* helpers.vhdl:221:43  */
  assign n31464_o = n31449_o[4];
  /* helpers.vhdl:221:43  */
  assign n31466_o = n31449_o[5];
  /* helpers.vhdl:221:43  */
  assign n31468_o = n31449_o[6];
  /* helpers.vhdl:221:43  */
  assign n31470_o = n31449_o[7];
  /* helpers.vhdl:221:43  */
  assign n31472_o = n31449_o[8];
  /* helpers.vhdl:221:43  */
  assign n31474_o = n31449_o[9];
  /* helpers.vhdl:221:43  */
  assign n31476_o = n31449_o[10];
  /* helpers.vhdl:221:43  */
  assign n31478_o = n31449_o[11];
  /* helpers.vhdl:221:43  */
  assign n31480_o = n31449_o[12];
  /* helpers.vhdl:221:43  */
  assign n31482_o = n31449_o[13];
  /* helpers.vhdl:221:43  */
  assign n31484_o = n31449_o[14];
  /* helpers.vhdl:221:43  */
  assign n31486_o = n31449_o[15];
  /* helpers.vhdl:221:43  */
  assign n31488_o = n31449_o[16];
  /* helpers.vhdl:221:43  */
  assign n31490_o = n31449_o[17];
  /* helpers.vhdl:221:43  */
  assign n31492_o = n31449_o[18];
  /* helpers.vhdl:221:43  */
  assign n31494_o = n31449_o[19];
  /* helpers.vhdl:221:43  */
  assign n31496_o = n31449_o[20];
  /* helpers.vhdl:221:43  */
  assign n31498_o = n31449_o[21];
  /* helpers.vhdl:221:43  */
  assign n31500_o = n31449_o[22];
  /* helpers.vhdl:221:43  */
  assign n31502_o = n31449_o[23];
  /* helpers.vhdl:221:43  */
  assign n31504_o = n31449_o[24];
  /* helpers.vhdl:221:43  */
  assign n31506_o = n31449_o[25];
  /* helpers.vhdl:221:43  */
  assign n31508_o = n31449_o[26];
  /* helpers.vhdl:221:43  */
  assign n31510_o = n31449_o[27];
  /* helpers.vhdl:221:43  */
  assign n31512_o = n31449_o[28];
  /* helpers.vhdl:221:43  */
  assign n31514_o = n31449_o[29];
  /* helpers.vhdl:221:43  */
  assign n31516_o = n31449_o[30];
  /* helpers.vhdl:221:43  */
  assign n31518_o = n31449_o[31];
  assign n31519_o = {n31455_o, n31458_o, n31460_o, n31462_o, n31464_o, n31466_o, n31468_o, n31470_o, n31472_o, n31474_o, n31476_o, n31478_o, n31480_o, n31482_o, n31484_o, n31486_o, n31488_o, n31490_o, n31492_o, n31494_o, n31496_o, n31498_o, n31500_o, n31502_o, n31504_o, n31506_o, n31508_o, n31510_o, n31512_o, n31514_o, n31516_o, n31518_o};
  /* countbits.vhdl:72:39  */
  assign n31520_o = rs[31:0];
  /* countbits.vhdl:69:13  */
  assign n31521_o = n31447_o ? n31519_o : n31520_o;
  assign n31522_o = {32'b11111111111111111111111111111111, n31521_o};
  /* countbits.vhdl:61:9  */
  assign n31523_o = n31308_o ? n31445_o : n31522_o;
  /* countbits.vhdl:76:49  */
  assign n31524_o = ~inp;
  /* countbits.vhdl:76:47  */
  assign n31526_o = {1'b0, n31524_o};
  /* countbits.vhdl:76:58  */
  assign n31528_o = n31526_o + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  /* countbits.vhdl:79:22  */
  assign n31529_o = sum_r[63:0];
  /* countbits.vhdl:79:36  */
  assign n31530_o = n31529_o | inp_r;
  /* helpers.vhdl:266:29  */
  assign n31540_o = \edge [1];
  /* helpers.vhdl:266:55  */
  assign n31541_o = \edge [0];
  /* helpers.vhdl:266:50  */
  assign n31542_o = ~n31541_o;
  /* helpers.vhdl:266:46  */
  assign n31543_o = n31540_o & n31542_o;
  /* helpers.vhdl:266:24  */
  assign n31545_o = 1'b0 | n31543_o;
  /* helpers.vhdl:266:29  */
  assign n31547_o = \edge [3];
  /* helpers.vhdl:266:55  */
  assign n31548_o = \edge [2];
  /* helpers.vhdl:266:50  */
  assign n31549_o = ~n31548_o;
  /* helpers.vhdl:266:46  */
  assign n31550_o = n31547_o & n31549_o;
  /* helpers.vhdl:266:24  */
  assign n31551_o = n31545_o | n31550_o;
  /* helpers.vhdl:266:29  */
  assign n31552_o = \edge [5];
  /* helpers.vhdl:266:55  */
  assign n31553_o = \edge [4];
  /* helpers.vhdl:266:50  */
  assign n31554_o = ~n31553_o;
  /* helpers.vhdl:266:46  */
  assign n31555_o = n31552_o & n31554_o;
  /* helpers.vhdl:266:24  */
  assign n31556_o = n31551_o | n31555_o;
  /* helpers.vhdl:266:29  */
  assign n31557_o = \edge [7];
  /* helpers.vhdl:266:55  */
  assign n31558_o = \edge [6];
  /* helpers.vhdl:266:50  */
  assign n31559_o = ~n31558_o;
  /* helpers.vhdl:266:46  */
  assign n31560_o = n31557_o & n31559_o;
  /* helpers.vhdl:266:24  */
  assign n31561_o = n31556_o | n31560_o;
  /* helpers.vhdl:266:29  */
  assign n31562_o = \edge [9];
  /* helpers.vhdl:266:55  */
  assign n31563_o = \edge [8];
  /* helpers.vhdl:266:50  */
  assign n31564_o = ~n31563_o;
  /* helpers.vhdl:266:46  */
  assign n31565_o = n31562_o & n31564_o;
  /* helpers.vhdl:266:24  */
  assign n31566_o = n31561_o | n31565_o;
  /* helpers.vhdl:266:29  */
  assign n31567_o = \edge [11];
  /* helpers.vhdl:266:55  */
  assign n31568_o = \edge [10];
  /* helpers.vhdl:266:50  */
  assign n31569_o = ~n31568_o;
  /* helpers.vhdl:266:46  */
  assign n31570_o = n31567_o & n31569_o;
  /* helpers.vhdl:266:24  */
  assign n31571_o = n31566_o | n31570_o;
  /* helpers.vhdl:266:29  */
  assign n31572_o = \edge [13];
  /* helpers.vhdl:266:55  */
  assign n31573_o = \edge [12];
  /* helpers.vhdl:266:50  */
  assign n31574_o = ~n31573_o;
  /* helpers.vhdl:266:46  */
  assign n31575_o = n31572_o & n31574_o;
  /* helpers.vhdl:266:24  */
  assign n31576_o = n31571_o | n31575_o;
  /* helpers.vhdl:266:29  */
  assign n31577_o = \edge [15];
  /* helpers.vhdl:266:55  */
  assign n31578_o = \edge [14];
  /* helpers.vhdl:266:50  */
  assign n31579_o = ~n31578_o;
  /* helpers.vhdl:266:46  */
  assign n31580_o = n31577_o & n31579_o;
  /* helpers.vhdl:266:24  */
  assign n31581_o = n31576_o | n31580_o;
  /* helpers.vhdl:266:29  */
  assign n31582_o = \edge [17];
  /* helpers.vhdl:266:55  */
  assign n31583_o = \edge [16];
  /* helpers.vhdl:266:50  */
  assign n31584_o = ~n31583_o;
  /* helpers.vhdl:266:46  */
  assign n31585_o = n31582_o & n31584_o;
  /* helpers.vhdl:266:24  */
  assign n31586_o = n31581_o | n31585_o;
  /* helpers.vhdl:266:29  */
  assign n31587_o = \edge [19];
  /* helpers.vhdl:266:55  */
  assign n31588_o = \edge [18];
  /* helpers.vhdl:266:50  */
  assign n31589_o = ~n31588_o;
  /* helpers.vhdl:266:46  */
  assign n31590_o = n31587_o & n31589_o;
  /* helpers.vhdl:266:24  */
  assign n31591_o = n31586_o | n31590_o;
  /* helpers.vhdl:266:29  */
  assign n31592_o = \edge [21];
  /* helpers.vhdl:266:55  */
  assign n31593_o = \edge [20];
  /* helpers.vhdl:266:50  */
  assign n31594_o = ~n31593_o;
  /* helpers.vhdl:266:46  */
  assign n31595_o = n31592_o & n31594_o;
  /* helpers.vhdl:266:24  */
  assign n31596_o = n31591_o | n31595_o;
  /* helpers.vhdl:266:29  */
  assign n31597_o = \edge [23];
  /* helpers.vhdl:266:55  */
  assign n31598_o = \edge [22];
  /* helpers.vhdl:266:50  */
  assign n31599_o = ~n31598_o;
  /* helpers.vhdl:266:46  */
  assign n31600_o = n31597_o & n31599_o;
  /* helpers.vhdl:266:24  */
  assign n31601_o = n31596_o | n31600_o;
  /* helpers.vhdl:266:29  */
  assign n31602_o = \edge [25];
  /* helpers.vhdl:266:55  */
  assign n31603_o = \edge [24];
  /* helpers.vhdl:266:50  */
  assign n31604_o = ~n31603_o;
  /* helpers.vhdl:266:46  */
  assign n31605_o = n31602_o & n31604_o;
  /* helpers.vhdl:266:24  */
  assign n31606_o = n31601_o | n31605_o;
  /* helpers.vhdl:266:29  */
  assign n31607_o = \edge [27];
  /* helpers.vhdl:266:55  */
  assign n31608_o = \edge [26];
  /* helpers.vhdl:266:50  */
  assign n31609_o = ~n31608_o;
  /* helpers.vhdl:266:46  */
  assign n31610_o = n31607_o & n31609_o;
  /* helpers.vhdl:266:24  */
  assign n31611_o = n31606_o | n31610_o;
  /* helpers.vhdl:266:29  */
  assign n31612_o = \edge [29];
  /* helpers.vhdl:266:55  */
  assign n31613_o = \edge [28];
  /* helpers.vhdl:266:50  */
  assign n31614_o = ~n31613_o;
  /* helpers.vhdl:266:46  */
  assign n31615_o = n31612_o & n31614_o;
  /* helpers.vhdl:266:24  */
  assign n31616_o = n31611_o | n31615_o;
  /* helpers.vhdl:266:29  */
  assign n31617_o = \edge [31];
  /* helpers.vhdl:266:55  */
  assign n31618_o = \edge [30];
  /* helpers.vhdl:266:50  */
  assign n31619_o = ~n31618_o;
  /* helpers.vhdl:266:46  */
  assign n31620_o = n31617_o & n31619_o;
  /* helpers.vhdl:266:24  */
  assign n31621_o = n31616_o | n31620_o;
  /* helpers.vhdl:266:29  */
  assign n31622_o = \edge [33];
  /* helpers.vhdl:266:55  */
  assign n31623_o = \edge [32];
  /* helpers.vhdl:266:50  */
  assign n31624_o = ~n31623_o;
  /* helpers.vhdl:266:46  */
  assign n31625_o = n31622_o & n31624_o;
  /* helpers.vhdl:266:24  */
  assign n31626_o = n31621_o | n31625_o;
  /* helpers.vhdl:266:29  */
  assign n31627_o = \edge [35];
  /* helpers.vhdl:266:55  */
  assign n31628_o = \edge [34];
  /* helpers.vhdl:266:50  */
  assign n31629_o = ~n31628_o;
  /* helpers.vhdl:266:46  */
  assign n31630_o = n31627_o & n31629_o;
  /* helpers.vhdl:266:24  */
  assign n31631_o = n31626_o | n31630_o;
  /* helpers.vhdl:266:29  */
  assign n31632_o = \edge [37];
  /* helpers.vhdl:266:55  */
  assign n31633_o = \edge [36];
  /* helpers.vhdl:266:50  */
  assign n31634_o = ~n31633_o;
  /* helpers.vhdl:266:46  */
  assign n31635_o = n31632_o & n31634_o;
  /* helpers.vhdl:266:24  */
  assign n31636_o = n31631_o | n31635_o;
  /* helpers.vhdl:266:29  */
  assign n31637_o = \edge [39];
  /* helpers.vhdl:266:55  */
  assign n31638_o = \edge [38];
  /* helpers.vhdl:266:50  */
  assign n31639_o = ~n31638_o;
  /* helpers.vhdl:266:46  */
  assign n31640_o = n31637_o & n31639_o;
  /* helpers.vhdl:266:24  */
  assign n31641_o = n31636_o | n31640_o;
  /* helpers.vhdl:266:29  */
  assign n31642_o = \edge [41];
  /* helpers.vhdl:266:55  */
  assign n31643_o = \edge [40];
  /* helpers.vhdl:266:50  */
  assign n31644_o = ~n31643_o;
  /* helpers.vhdl:266:46  */
  assign n31645_o = n31642_o & n31644_o;
  /* helpers.vhdl:266:24  */
  assign n31646_o = n31641_o | n31645_o;
  /* helpers.vhdl:266:29  */
  assign n31647_o = \edge [43];
  /* helpers.vhdl:266:55  */
  assign n31648_o = \edge [42];
  /* helpers.vhdl:266:50  */
  assign n31649_o = ~n31648_o;
  /* helpers.vhdl:266:46  */
  assign n31650_o = n31647_o & n31649_o;
  /* helpers.vhdl:266:24  */
  assign n31651_o = n31646_o | n31650_o;
  /* helpers.vhdl:266:29  */
  assign n31652_o = \edge [45];
  /* helpers.vhdl:266:55  */
  assign n31653_o = \edge [44];
  /* helpers.vhdl:266:50  */
  assign n31654_o = ~n31653_o;
  /* helpers.vhdl:266:46  */
  assign n31655_o = n31652_o & n31654_o;
  /* helpers.vhdl:266:24  */
  assign n31656_o = n31651_o | n31655_o;
  /* helpers.vhdl:266:29  */
  assign n31657_o = \edge [47];
  /* helpers.vhdl:266:55  */
  assign n31658_o = \edge [46];
  /* helpers.vhdl:266:50  */
  assign n31659_o = ~n31658_o;
  /* helpers.vhdl:266:46  */
  assign n31660_o = n31657_o & n31659_o;
  /* helpers.vhdl:266:24  */
  assign n31661_o = n31656_o | n31660_o;
  /* helpers.vhdl:266:29  */
  assign n31662_o = \edge [49];
  /* helpers.vhdl:266:55  */
  assign n31663_o = \edge [48];
  /* helpers.vhdl:266:50  */
  assign n31664_o = ~n31663_o;
  /* helpers.vhdl:266:46  */
  assign n31665_o = n31662_o & n31664_o;
  /* helpers.vhdl:266:24  */
  assign n31666_o = n31661_o | n31665_o;
  /* helpers.vhdl:266:29  */
  assign n31667_o = \edge [51];
  /* helpers.vhdl:266:55  */
  assign n31668_o = \edge [50];
  /* helpers.vhdl:266:50  */
  assign n31669_o = ~n31668_o;
  /* helpers.vhdl:266:46  */
  assign n31670_o = n31667_o & n31669_o;
  /* helpers.vhdl:266:24  */
  assign n31671_o = n31666_o | n31670_o;
  /* helpers.vhdl:266:29  */
  assign n31672_o = \edge [53];
  /* helpers.vhdl:266:55  */
  assign n31673_o = \edge [52];
  /* helpers.vhdl:266:50  */
  assign n31674_o = ~n31673_o;
  /* helpers.vhdl:266:46  */
  assign n31675_o = n31672_o & n31674_o;
  /* helpers.vhdl:266:24  */
  assign n31676_o = n31671_o | n31675_o;
  /* helpers.vhdl:266:29  */
  assign n31677_o = \edge [55];
  /* helpers.vhdl:266:55  */
  assign n31678_o = \edge [54];
  /* helpers.vhdl:266:50  */
  assign n31679_o = ~n31678_o;
  /* helpers.vhdl:266:46  */
  assign n31680_o = n31677_o & n31679_o;
  /* helpers.vhdl:266:24  */
  assign n31681_o = n31676_o | n31680_o;
  /* helpers.vhdl:266:29  */
  assign n31682_o = \edge [57];
  /* helpers.vhdl:266:55  */
  assign n31683_o = \edge [56];
  /* helpers.vhdl:266:50  */
  assign n31684_o = ~n31683_o;
  /* helpers.vhdl:266:46  */
  assign n31685_o = n31682_o & n31684_o;
  /* helpers.vhdl:266:24  */
  assign n31686_o = n31681_o | n31685_o;
  /* helpers.vhdl:266:29  */
  assign n31687_o = \edge [59];
  /* helpers.vhdl:266:55  */
  assign n31688_o = \edge [58];
  /* helpers.vhdl:266:50  */
  assign n31689_o = ~n31688_o;
  /* helpers.vhdl:266:46  */
  assign n31690_o = n31687_o & n31689_o;
  /* helpers.vhdl:266:24  */
  assign n31691_o = n31686_o | n31690_o;
  /* helpers.vhdl:266:29  */
  assign n31692_o = \edge [61];
  /* helpers.vhdl:266:55  */
  assign n31693_o = \edge [60];
  /* helpers.vhdl:266:50  */
  assign n31694_o = ~n31693_o;
  /* helpers.vhdl:266:46  */
  assign n31695_o = n31692_o & n31694_o;
  /* helpers.vhdl:266:24  */
  assign n31696_o = n31691_o | n31695_o;
  /* helpers.vhdl:266:29  */
  assign n31697_o = \edge [63];
  /* helpers.vhdl:266:55  */
  assign n31698_o = \edge [62];
  /* helpers.vhdl:266:50  */
  assign n31699_o = ~n31698_o;
  /* helpers.vhdl:266:46  */
  assign n31700_o = n31697_o & n31699_o;
  /* helpers.vhdl:266:24  */
  assign n31701_o = n31696_o | n31700_o;
  /* helpers.vhdl:266:29  */
  assign n31704_o = \edge [3];
  /* helpers.vhdl:266:55  */
  assign n31705_o = \edge [1];
  /* helpers.vhdl:266:50  */
  assign n31706_o = ~n31705_o;
  /* helpers.vhdl:266:46  */
  assign n31707_o = n31704_o & n31706_o;
  /* helpers.vhdl:266:24  */
  assign n31709_o = 1'b0 | n31707_o;
  /* helpers.vhdl:266:29  */
  assign n31711_o = \edge [7];
  /* helpers.vhdl:266:55  */
  assign n31712_o = \edge [5];
  /* helpers.vhdl:266:50  */
  assign n31713_o = ~n31712_o;
  /* helpers.vhdl:266:46  */
  assign n31714_o = n31711_o & n31713_o;
  /* helpers.vhdl:266:24  */
  assign n31715_o = n31709_o | n31714_o;
  /* helpers.vhdl:266:29  */
  assign n31716_o = \edge [11];
  /* helpers.vhdl:266:55  */
  assign n31717_o = \edge [9];
  /* helpers.vhdl:266:50  */
  assign n31718_o = ~n31717_o;
  /* helpers.vhdl:266:46  */
  assign n31719_o = n31716_o & n31718_o;
  /* helpers.vhdl:266:24  */
  assign n31720_o = n31715_o | n31719_o;
  /* helpers.vhdl:266:29  */
  assign n31721_o = \edge [15];
  /* helpers.vhdl:266:55  */
  assign n31722_o = \edge [13];
  /* helpers.vhdl:266:50  */
  assign n31723_o = ~n31722_o;
  /* helpers.vhdl:266:46  */
  assign n31724_o = n31721_o & n31723_o;
  /* helpers.vhdl:266:24  */
  assign n31725_o = n31720_o | n31724_o;
  /* helpers.vhdl:266:29  */
  assign n31726_o = \edge [19];
  /* helpers.vhdl:266:55  */
  assign n31727_o = \edge [17];
  /* helpers.vhdl:266:50  */
  assign n31728_o = ~n31727_o;
  /* helpers.vhdl:266:46  */
  assign n31729_o = n31726_o & n31728_o;
  /* helpers.vhdl:266:24  */
  assign n31730_o = n31725_o | n31729_o;
  /* helpers.vhdl:266:29  */
  assign n31731_o = \edge [23];
  /* helpers.vhdl:266:55  */
  assign n31732_o = \edge [21];
  /* helpers.vhdl:266:50  */
  assign n31733_o = ~n31732_o;
  /* helpers.vhdl:266:46  */
  assign n31734_o = n31731_o & n31733_o;
  /* helpers.vhdl:266:24  */
  assign n31735_o = n31730_o | n31734_o;
  /* helpers.vhdl:266:29  */
  assign n31736_o = \edge [27];
  /* helpers.vhdl:266:55  */
  assign n31737_o = \edge [25];
  /* helpers.vhdl:266:50  */
  assign n31738_o = ~n31737_o;
  /* helpers.vhdl:266:46  */
  assign n31739_o = n31736_o & n31738_o;
  /* helpers.vhdl:266:24  */
  assign n31740_o = n31735_o | n31739_o;
  /* helpers.vhdl:266:29  */
  assign n31741_o = \edge [31];
  /* helpers.vhdl:266:55  */
  assign n31742_o = \edge [29];
  /* helpers.vhdl:266:50  */
  assign n31743_o = ~n31742_o;
  /* helpers.vhdl:266:46  */
  assign n31744_o = n31741_o & n31743_o;
  /* helpers.vhdl:266:24  */
  assign n31745_o = n31740_o | n31744_o;
  /* helpers.vhdl:266:29  */
  assign n31746_o = \edge [35];
  /* helpers.vhdl:266:55  */
  assign n31747_o = \edge [33];
  /* helpers.vhdl:266:50  */
  assign n31748_o = ~n31747_o;
  /* helpers.vhdl:266:46  */
  assign n31749_o = n31746_o & n31748_o;
  /* helpers.vhdl:266:24  */
  assign n31750_o = n31745_o | n31749_o;
  /* helpers.vhdl:266:29  */
  assign n31751_o = \edge [39];
  /* helpers.vhdl:266:55  */
  assign n31752_o = \edge [37];
  /* helpers.vhdl:266:50  */
  assign n31753_o = ~n31752_o;
  /* helpers.vhdl:266:46  */
  assign n31754_o = n31751_o & n31753_o;
  /* helpers.vhdl:266:24  */
  assign n31755_o = n31750_o | n31754_o;
  /* helpers.vhdl:266:29  */
  assign n31756_o = \edge [43];
  /* helpers.vhdl:266:55  */
  assign n31757_o = \edge [41];
  /* helpers.vhdl:266:50  */
  assign n31758_o = ~n31757_o;
  /* helpers.vhdl:266:46  */
  assign n31759_o = n31756_o & n31758_o;
  /* helpers.vhdl:266:24  */
  assign n31760_o = n31755_o | n31759_o;
  /* helpers.vhdl:266:29  */
  assign n31761_o = \edge [47];
  /* helpers.vhdl:266:55  */
  assign n31762_o = \edge [45];
  /* helpers.vhdl:266:50  */
  assign n31763_o = ~n31762_o;
  /* helpers.vhdl:266:46  */
  assign n31764_o = n31761_o & n31763_o;
  /* helpers.vhdl:266:24  */
  assign n31765_o = n31760_o | n31764_o;
  /* helpers.vhdl:266:29  */
  assign n31766_o = \edge [51];
  /* helpers.vhdl:266:55  */
  assign n31767_o = \edge [49];
  /* helpers.vhdl:266:50  */
  assign n31768_o = ~n31767_o;
  /* helpers.vhdl:266:46  */
  assign n31769_o = n31766_o & n31768_o;
  /* helpers.vhdl:266:24  */
  assign n31770_o = n31765_o | n31769_o;
  /* helpers.vhdl:266:29  */
  assign n31771_o = \edge [55];
  /* helpers.vhdl:266:55  */
  assign n31772_o = \edge [53];
  /* helpers.vhdl:266:50  */
  assign n31773_o = ~n31772_o;
  /* helpers.vhdl:266:46  */
  assign n31774_o = n31771_o & n31773_o;
  /* helpers.vhdl:266:24  */
  assign n31775_o = n31770_o | n31774_o;
  /* helpers.vhdl:266:29  */
  assign n31776_o = \edge [59];
  /* helpers.vhdl:266:55  */
  assign n31777_o = \edge [57];
  /* helpers.vhdl:266:50  */
  assign n31778_o = ~n31777_o;
  /* helpers.vhdl:266:46  */
  assign n31779_o = n31776_o & n31778_o;
  /* helpers.vhdl:266:24  */
  assign n31780_o = n31775_o | n31779_o;
  /* helpers.vhdl:266:29  */
  assign n31781_o = \edge [63];
  /* helpers.vhdl:266:55  */
  assign n31782_o = \edge [61];
  /* helpers.vhdl:266:50  */
  assign n31783_o = ~n31782_o;
  /* helpers.vhdl:266:46  */
  assign n31784_o = n31781_o & n31783_o;
  /* helpers.vhdl:266:24  */
  assign n31785_o = n31780_o | n31784_o;
  /* helpers.vhdl:266:29  */
  assign n31787_o = \edge [7];
  /* helpers.vhdl:266:55  */
  assign n31788_o = \edge [3];
  /* helpers.vhdl:266:50  */
  assign n31789_o = ~n31788_o;
  /* helpers.vhdl:266:46  */
  assign n31790_o = n31787_o & n31789_o;
  /* helpers.vhdl:266:24  */
  assign n31792_o = 1'b0 | n31790_o;
  /* helpers.vhdl:266:29  */
  assign n31794_o = \edge [15];
  /* helpers.vhdl:266:55  */
  assign n31795_o = \edge [11];
  /* helpers.vhdl:266:50  */
  assign n31796_o = ~n31795_o;
  /* helpers.vhdl:266:46  */
  assign n31797_o = n31794_o & n31796_o;
  /* helpers.vhdl:266:24  */
  assign n31798_o = n31792_o | n31797_o;
  /* helpers.vhdl:266:29  */
  assign n31799_o = \edge [23];
  /* helpers.vhdl:266:55  */
  assign n31800_o = \edge [19];
  /* helpers.vhdl:266:50  */
  assign n31801_o = ~n31800_o;
  /* helpers.vhdl:266:46  */
  assign n31802_o = n31799_o & n31801_o;
  /* helpers.vhdl:266:24  */
  assign n31803_o = n31798_o | n31802_o;
  /* helpers.vhdl:266:29  */
  assign n31804_o = \edge [31];
  /* helpers.vhdl:266:55  */
  assign n31805_o = \edge [27];
  /* helpers.vhdl:266:50  */
  assign n31806_o = ~n31805_o;
  /* helpers.vhdl:266:46  */
  assign n31807_o = n31804_o & n31806_o;
  /* helpers.vhdl:266:24  */
  assign n31808_o = n31803_o | n31807_o;
  /* helpers.vhdl:266:29  */
  assign n31809_o = \edge [39];
  /* helpers.vhdl:266:55  */
  assign n31810_o = \edge [35];
  /* helpers.vhdl:266:50  */
  assign n31811_o = ~n31810_o;
  /* helpers.vhdl:266:46  */
  assign n31812_o = n31809_o & n31811_o;
  /* helpers.vhdl:266:24  */
  assign n31813_o = n31808_o | n31812_o;
  /* helpers.vhdl:266:29  */
  assign n31814_o = \edge [47];
  /* helpers.vhdl:266:55  */
  assign n31815_o = \edge [43];
  /* helpers.vhdl:266:50  */
  assign n31816_o = ~n31815_o;
  /* helpers.vhdl:266:46  */
  assign n31817_o = n31814_o & n31816_o;
  /* helpers.vhdl:266:24  */
  assign n31818_o = n31813_o | n31817_o;
  /* helpers.vhdl:266:29  */
  assign n31819_o = \edge [55];
  /* helpers.vhdl:266:55  */
  assign n31820_o = \edge [51];
  /* helpers.vhdl:266:50  */
  assign n31821_o = ~n31820_o;
  /* helpers.vhdl:266:46  */
  assign n31822_o = n31819_o & n31821_o;
  /* helpers.vhdl:266:24  */
  assign n31823_o = n31818_o | n31822_o;
  /* helpers.vhdl:266:29  */
  assign n31824_o = \edge [63];
  /* helpers.vhdl:266:55  */
  assign n31825_o = \edge [59];
  /* helpers.vhdl:266:50  */
  assign n31826_o = ~n31825_o;
  /* helpers.vhdl:266:46  */
  assign n31827_o = n31824_o & n31826_o;
  /* helpers.vhdl:266:24  */
  assign n31828_o = n31823_o | n31827_o;
  /* helpers.vhdl:266:29  */
  assign n31830_o = \edge [15];
  /* helpers.vhdl:266:55  */
  assign n31831_o = \edge [7];
  /* helpers.vhdl:266:50  */
  assign n31832_o = ~n31831_o;
  /* helpers.vhdl:266:46  */
  assign n31833_o = n31830_o & n31832_o;
  /* helpers.vhdl:266:24  */
  assign n31835_o = 1'b0 | n31833_o;
  /* helpers.vhdl:266:29  */
  assign n31837_o = \edge [31];
  /* helpers.vhdl:266:55  */
  assign n31838_o = \edge [23];
  /* helpers.vhdl:266:50  */
  assign n31839_o = ~n31838_o;
  /* helpers.vhdl:266:46  */
  assign n31840_o = n31837_o & n31839_o;
  /* helpers.vhdl:266:24  */
  assign n31841_o = n31835_o | n31840_o;
  /* helpers.vhdl:266:29  */
  assign n31842_o = \edge [47];
  /* helpers.vhdl:266:55  */
  assign n31843_o = \edge [39];
  /* helpers.vhdl:266:50  */
  assign n31844_o = ~n31843_o;
  /* helpers.vhdl:266:46  */
  assign n31845_o = n31842_o & n31844_o;
  /* helpers.vhdl:266:24  */
  assign n31846_o = n31841_o | n31845_o;
  /* helpers.vhdl:266:29  */
  assign n31847_o = \edge [63];
  /* helpers.vhdl:266:55  */
  assign n31848_o = \edge [55];
  /* helpers.vhdl:266:50  */
  assign n31849_o = ~n31848_o;
  /* helpers.vhdl:266:46  */
  assign n31850_o = n31847_o & n31849_o;
  /* helpers.vhdl:266:24  */
  assign n31851_o = n31846_o | n31850_o;
  /* helpers.vhdl:266:29  */
  assign n31853_o = \edge [31];
  /* helpers.vhdl:266:55  */
  assign n31854_o = \edge [15];
  /* helpers.vhdl:266:50  */
  assign n31855_o = ~n31854_o;
  /* helpers.vhdl:266:46  */
  assign n31856_o = n31853_o & n31855_o;
  /* helpers.vhdl:266:24  */
  assign n31858_o = 1'b0 | n31856_o;
  /* helpers.vhdl:266:29  */
  assign n31860_o = \edge [63];
  /* helpers.vhdl:266:55  */
  assign n31861_o = \edge [47];
  /* helpers.vhdl:266:50  */
  assign n31862_o = ~n31861_o;
  /* helpers.vhdl:266:46  */
  assign n31863_o = n31860_o & n31862_o;
  /* helpers.vhdl:266:24  */
  assign n31864_o = n31858_o | n31863_o;
  /* helpers.vhdl:266:29  */
  assign n31866_o = \edge [63];
  /* helpers.vhdl:266:55  */
  assign n31867_o = \edge [31];
  /* helpers.vhdl:266:50  */
  assign n31868_o = ~n31867_o;
  /* helpers.vhdl:266:46  */
  assign n31869_o = n31866_o & n31868_o;
  /* helpers.vhdl:266:24  */
  assign n31871_o = 1'b0 | n31869_o;
  assign n31873_o = {n31871_o, n31864_o, n31851_o, n31828_o, n31785_o, n31701_o};
  /* countbits.vhdl:81:24  */
  assign n31874_o = sum_r[63:0];
  /* countbits.vhdl:81:38  */
  assign n31875_o = n31874_o & inp_r;
  /* helpers.vhdl:244:36  */
  assign n31885_o = onehot[1];
  /* helpers.vhdl:244:32  */
  assign n31886_o = |(n31885_o);
  /* helpers.vhdl:244:28  */
  assign n31888_o = 1'b0 | n31886_o;
  /* helpers.vhdl:244:36  */
  assign n31890_o = onehot[3];
  /* helpers.vhdl:244:32  */
  assign n31891_o = |(n31890_o);
  /* helpers.vhdl:244:28  */
  assign n31892_o = n31888_o | n31891_o;
  /* helpers.vhdl:244:36  */
  assign n31893_o = onehot[5];
  /* helpers.vhdl:244:32  */
  assign n31894_o = |(n31893_o);
  /* helpers.vhdl:244:28  */
  assign n31895_o = n31892_o | n31894_o;
  /* helpers.vhdl:244:36  */
  assign n31896_o = onehot[7];
  /* helpers.vhdl:244:32  */
  assign n31897_o = |(n31896_o);
  /* helpers.vhdl:244:28  */
  assign n31898_o = n31895_o | n31897_o;
  /* helpers.vhdl:244:36  */
  assign n31899_o = onehot[9];
  /* helpers.vhdl:244:32  */
  assign n31900_o = |(n31899_o);
  /* helpers.vhdl:244:28  */
  assign n31901_o = n31898_o | n31900_o;
  /* helpers.vhdl:244:36  */
  assign n31902_o = onehot[11];
  /* helpers.vhdl:244:32  */
  assign n31903_o = |(n31902_o);
  /* helpers.vhdl:244:28  */
  assign n31904_o = n31901_o | n31903_o;
  /* helpers.vhdl:244:36  */
  assign n31905_o = onehot[13];
  /* helpers.vhdl:244:32  */
  assign n31906_o = |(n31905_o);
  /* helpers.vhdl:244:28  */
  assign n31907_o = n31904_o | n31906_o;
  /* helpers.vhdl:244:36  */
  assign n31908_o = onehot[15];
  /* helpers.vhdl:244:32  */
  assign n31909_o = |(n31908_o);
  /* helpers.vhdl:244:28  */
  assign n31910_o = n31907_o | n31909_o;
  /* helpers.vhdl:244:36  */
  assign n31911_o = onehot[17];
  /* helpers.vhdl:244:32  */
  assign n31912_o = |(n31911_o);
  /* helpers.vhdl:244:28  */
  assign n31913_o = n31910_o | n31912_o;
  /* helpers.vhdl:244:36  */
  assign n31914_o = onehot[19];
  /* helpers.vhdl:244:32  */
  assign n31915_o = |(n31914_o);
  /* helpers.vhdl:244:28  */
  assign n31916_o = n31913_o | n31915_o;
  /* helpers.vhdl:244:36  */
  assign n31917_o = onehot[21];
  /* helpers.vhdl:244:32  */
  assign n31918_o = |(n31917_o);
  /* helpers.vhdl:244:28  */
  assign n31919_o = n31916_o | n31918_o;
  /* helpers.vhdl:244:36  */
  assign n31920_o = onehot[23];
  /* helpers.vhdl:244:32  */
  assign n31921_o = |(n31920_o);
  /* helpers.vhdl:244:28  */
  assign n31922_o = n31919_o | n31921_o;
  /* helpers.vhdl:244:36  */
  assign n31923_o = onehot[25];
  /* helpers.vhdl:244:32  */
  assign n31924_o = |(n31923_o);
  /* helpers.vhdl:244:28  */
  assign n31925_o = n31922_o | n31924_o;
  /* helpers.vhdl:244:36  */
  assign n31926_o = onehot[27];
  /* helpers.vhdl:244:32  */
  assign n31927_o = |(n31926_o);
  /* helpers.vhdl:244:28  */
  assign n31928_o = n31925_o | n31927_o;
  /* helpers.vhdl:244:36  */
  assign n31929_o = onehot[29];
  /* helpers.vhdl:244:32  */
  assign n31930_o = |(n31929_o);
  /* helpers.vhdl:244:28  */
  assign n31931_o = n31928_o | n31930_o;
  /* helpers.vhdl:244:36  */
  assign n31932_o = onehot[31];
  /* helpers.vhdl:244:32  */
  assign n31933_o = |(n31932_o);
  /* helpers.vhdl:244:28  */
  assign n31934_o = n31931_o | n31933_o;
  /* helpers.vhdl:244:36  */
  assign n31935_o = onehot[33];
  /* helpers.vhdl:244:32  */
  assign n31936_o = |(n31935_o);
  /* helpers.vhdl:244:28  */
  assign n31937_o = n31934_o | n31936_o;
  /* helpers.vhdl:244:36  */
  assign n31938_o = onehot[35];
  /* helpers.vhdl:244:32  */
  assign n31939_o = |(n31938_o);
  /* helpers.vhdl:244:28  */
  assign n31940_o = n31937_o | n31939_o;
  /* helpers.vhdl:244:36  */
  assign n31941_o = onehot[37];
  /* helpers.vhdl:244:32  */
  assign n31942_o = |(n31941_o);
  /* helpers.vhdl:244:28  */
  assign n31943_o = n31940_o | n31942_o;
  /* helpers.vhdl:244:36  */
  assign n31944_o = onehot[39];
  /* helpers.vhdl:244:32  */
  assign n31945_o = |(n31944_o);
  /* helpers.vhdl:244:28  */
  assign n31946_o = n31943_o | n31945_o;
  /* helpers.vhdl:244:36  */
  assign n31947_o = onehot[41];
  /* helpers.vhdl:244:32  */
  assign n31948_o = |(n31947_o);
  /* helpers.vhdl:244:28  */
  assign n31949_o = n31946_o | n31948_o;
  /* helpers.vhdl:244:36  */
  assign n31950_o = onehot[43];
  /* helpers.vhdl:244:32  */
  assign n31951_o = |(n31950_o);
  /* helpers.vhdl:244:28  */
  assign n31952_o = n31949_o | n31951_o;
  /* helpers.vhdl:244:36  */
  assign n31953_o = onehot[45];
  /* helpers.vhdl:244:32  */
  assign n31954_o = |(n31953_o);
  /* helpers.vhdl:244:28  */
  assign n31955_o = n31952_o | n31954_o;
  /* helpers.vhdl:244:36  */
  assign n31956_o = onehot[47];
  /* helpers.vhdl:244:32  */
  assign n31957_o = |(n31956_o);
  /* helpers.vhdl:244:28  */
  assign n31958_o = n31955_o | n31957_o;
  /* helpers.vhdl:244:36  */
  assign n31959_o = onehot[49];
  /* helpers.vhdl:244:32  */
  assign n31960_o = |(n31959_o);
  /* helpers.vhdl:244:28  */
  assign n31961_o = n31958_o | n31960_o;
  /* helpers.vhdl:244:36  */
  assign n31962_o = onehot[51];
  /* helpers.vhdl:244:32  */
  assign n31963_o = |(n31962_o);
  /* helpers.vhdl:244:28  */
  assign n31964_o = n31961_o | n31963_o;
  /* helpers.vhdl:244:36  */
  assign n31965_o = onehot[53];
  /* helpers.vhdl:244:32  */
  assign n31966_o = |(n31965_o);
  /* helpers.vhdl:244:28  */
  assign n31967_o = n31964_o | n31966_o;
  /* helpers.vhdl:244:36  */
  assign n31968_o = onehot[55];
  /* helpers.vhdl:244:32  */
  assign n31969_o = |(n31968_o);
  /* helpers.vhdl:244:28  */
  assign n31970_o = n31967_o | n31969_o;
  /* helpers.vhdl:244:36  */
  assign n31971_o = onehot[57];
  /* helpers.vhdl:244:32  */
  assign n31972_o = |(n31971_o);
  /* helpers.vhdl:244:28  */
  assign n31973_o = n31970_o | n31972_o;
  /* helpers.vhdl:244:36  */
  assign n31974_o = onehot[59];
  /* helpers.vhdl:244:32  */
  assign n31975_o = |(n31974_o);
  /* helpers.vhdl:244:28  */
  assign n31976_o = n31973_o | n31975_o;
  /* helpers.vhdl:244:36  */
  assign n31977_o = onehot[61];
  /* helpers.vhdl:244:32  */
  assign n31978_o = |(n31977_o);
  /* helpers.vhdl:244:28  */
  assign n31979_o = n31976_o | n31978_o;
  /* helpers.vhdl:244:36  */
  assign n31980_o = onehot[63];
  /* helpers.vhdl:244:32  */
  assign n31981_o = |(n31980_o);
  /* helpers.vhdl:244:28  */
  assign n31982_o = n31979_o | n31981_o;
  /* helpers.vhdl:244:36  */
  assign n31985_o = onehot[3:2];
  /* helpers.vhdl:244:32  */
  assign n31986_o = |(n31985_o);
  /* helpers.vhdl:244:28  */
  assign n31988_o = 1'b0 | n31986_o;
  /* helpers.vhdl:244:36  */
  assign n31990_o = onehot[7:6];
  /* helpers.vhdl:244:32  */
  assign n31991_o = |(n31990_o);
  /* helpers.vhdl:244:28  */
  assign n31992_o = n31988_o | n31991_o;
  /* helpers.vhdl:244:36  */
  assign n31993_o = onehot[11:10];
  /* helpers.vhdl:244:32  */
  assign n31994_o = |(n31993_o);
  /* helpers.vhdl:244:28  */
  assign n31995_o = n31992_o | n31994_o;
  /* helpers.vhdl:244:36  */
  assign n31996_o = onehot[15:14];
  /* helpers.vhdl:244:32  */
  assign n31997_o = |(n31996_o);
  /* helpers.vhdl:244:28  */
  assign n31998_o = n31995_o | n31997_o;
  /* helpers.vhdl:244:36  */
  assign n31999_o = onehot[19:18];
  /* helpers.vhdl:244:32  */
  assign n32000_o = |(n31999_o);
  /* helpers.vhdl:244:28  */
  assign n32001_o = n31998_o | n32000_o;
  /* helpers.vhdl:244:36  */
  assign n32002_o = onehot[23:22];
  /* helpers.vhdl:244:32  */
  assign n32003_o = |(n32002_o);
  /* helpers.vhdl:244:28  */
  assign n32004_o = n32001_o | n32003_o;
  /* helpers.vhdl:244:36  */
  assign n32005_o = onehot[27:26];
  /* helpers.vhdl:244:32  */
  assign n32006_o = |(n32005_o);
  /* helpers.vhdl:244:28  */
  assign n32007_o = n32004_o | n32006_o;
  /* helpers.vhdl:244:36  */
  assign n32008_o = onehot[31:30];
  /* helpers.vhdl:244:32  */
  assign n32009_o = |(n32008_o);
  /* helpers.vhdl:244:28  */
  assign n32010_o = n32007_o | n32009_o;
  /* helpers.vhdl:244:36  */
  assign n32011_o = onehot[35:34];
  /* helpers.vhdl:244:32  */
  assign n32012_o = |(n32011_o);
  /* helpers.vhdl:244:28  */
  assign n32013_o = n32010_o | n32012_o;
  /* helpers.vhdl:244:36  */
  assign n32014_o = onehot[39:38];
  /* helpers.vhdl:244:32  */
  assign n32015_o = |(n32014_o);
  /* helpers.vhdl:244:28  */
  assign n32016_o = n32013_o | n32015_o;
  /* helpers.vhdl:244:36  */
  assign n32017_o = onehot[43:42];
  /* helpers.vhdl:244:32  */
  assign n32018_o = |(n32017_o);
  /* helpers.vhdl:244:28  */
  assign n32019_o = n32016_o | n32018_o;
  /* helpers.vhdl:244:36  */
  assign n32020_o = onehot[47:46];
  /* helpers.vhdl:244:32  */
  assign n32021_o = |(n32020_o);
  /* helpers.vhdl:244:28  */
  assign n32022_o = n32019_o | n32021_o;
  /* helpers.vhdl:244:36  */
  assign n32023_o = onehot[51:50];
  /* helpers.vhdl:244:32  */
  assign n32024_o = |(n32023_o);
  /* helpers.vhdl:244:28  */
  assign n32025_o = n32022_o | n32024_o;
  /* helpers.vhdl:244:36  */
  assign n32026_o = onehot[55:54];
  /* helpers.vhdl:244:32  */
  assign n32027_o = |(n32026_o);
  /* helpers.vhdl:244:28  */
  assign n32028_o = n32025_o | n32027_o;
  /* helpers.vhdl:244:36  */
  assign n32029_o = onehot[59:58];
  /* helpers.vhdl:244:32  */
  assign n32030_o = |(n32029_o);
  /* helpers.vhdl:244:28  */
  assign n32031_o = n32028_o | n32030_o;
  /* helpers.vhdl:244:36  */
  assign n32032_o = onehot[63:62];
  /* helpers.vhdl:244:32  */
  assign n32033_o = |(n32032_o);
  /* helpers.vhdl:244:28  */
  assign n32034_o = n32031_o | n32033_o;
  /* helpers.vhdl:244:36  */
  assign n32036_o = onehot[7:4];
  /* helpers.vhdl:244:32  */
  assign n32037_o = |(n32036_o);
  /* helpers.vhdl:244:28  */
  assign n32039_o = 1'b0 | n32037_o;
  /* helpers.vhdl:244:36  */
  assign n32041_o = onehot[15:12];
  /* helpers.vhdl:244:32  */
  assign n32042_o = |(n32041_o);
  /* helpers.vhdl:244:28  */
  assign n32043_o = n32039_o | n32042_o;
  /* helpers.vhdl:244:36  */
  assign n32044_o = onehot[23:20];
  /* helpers.vhdl:244:32  */
  assign n32045_o = |(n32044_o);
  /* helpers.vhdl:244:28  */
  assign n32046_o = n32043_o | n32045_o;
  /* helpers.vhdl:244:36  */
  assign n32047_o = onehot[31:28];
  /* helpers.vhdl:244:32  */
  assign n32048_o = |(n32047_o);
  /* helpers.vhdl:244:28  */
  assign n32049_o = n32046_o | n32048_o;
  /* helpers.vhdl:244:36  */
  assign n32050_o = onehot[39:36];
  /* helpers.vhdl:244:32  */
  assign n32051_o = |(n32050_o);
  /* helpers.vhdl:244:28  */
  assign n32052_o = n32049_o | n32051_o;
  /* helpers.vhdl:244:36  */
  assign n32053_o = onehot[47:44];
  /* helpers.vhdl:244:32  */
  assign n32054_o = |(n32053_o);
  /* helpers.vhdl:244:28  */
  assign n32055_o = n32052_o | n32054_o;
  /* helpers.vhdl:244:36  */
  assign n32056_o = onehot[55:52];
  /* helpers.vhdl:244:32  */
  assign n32057_o = |(n32056_o);
  /* helpers.vhdl:244:28  */
  assign n32058_o = n32055_o | n32057_o;
  /* helpers.vhdl:244:36  */
  assign n32059_o = onehot[63:60];
  /* helpers.vhdl:244:32  */
  assign n32060_o = |(n32059_o);
  /* helpers.vhdl:244:28  */
  assign n32061_o = n32058_o | n32060_o;
  /* helpers.vhdl:244:36  */
  assign n32063_o = onehot[15:8];
  /* helpers.vhdl:244:32  */
  assign n32064_o = |(n32063_o);
  /* helpers.vhdl:244:28  */
  assign n32066_o = 1'b0 | n32064_o;
  /* helpers.vhdl:244:36  */
  assign n32068_o = onehot[31:24];
  /* helpers.vhdl:244:32  */
  assign n32069_o = |(n32068_o);
  /* helpers.vhdl:244:28  */
  assign n32070_o = n32066_o | n32069_o;
  /* helpers.vhdl:244:36  */
  assign n32071_o = onehot[47:40];
  /* helpers.vhdl:244:32  */
  assign n32072_o = |(n32071_o);
  /* helpers.vhdl:244:28  */
  assign n32073_o = n32070_o | n32072_o;
  /* helpers.vhdl:244:36  */
  assign n32074_o = onehot[63:56];
  /* helpers.vhdl:244:32  */
  assign n32075_o = |(n32074_o);
  /* helpers.vhdl:244:28  */
  assign n32076_o = n32073_o | n32075_o;
  /* helpers.vhdl:244:36  */
  assign n32078_o = onehot[31:16];
  /* helpers.vhdl:244:32  */
  assign n32079_o = |(n32078_o);
  /* helpers.vhdl:244:28  */
  assign n32081_o = 1'b0 | n32079_o;
  /* helpers.vhdl:244:36  */
  assign n32083_o = onehot[63:48];
  /* helpers.vhdl:244:32  */
  assign n32084_o = |(n32083_o);
  /* helpers.vhdl:244:28  */
  assign n32085_o = n32081_o | n32084_o;
  /* helpers.vhdl:244:36  */
  assign n32087_o = onehot[63:32];
  /* helpers.vhdl:244:32  */
  assign n32088_o = |(n32087_o);
  /* helpers.vhdl:244:28  */
  assign n32090_o = 1'b0 | n32088_o;
  assign n32092_o = {n32090_o, n32085_o, n32076_o, n32061_o, n32034_o, n31982_o};
  /* countbits.vhdl:83:39  */
  assign n32093_o = n31873_o[5:2];
  /* countbits.vhdl:84:39  */
  assign n32094_o = n32092_o[1:0];
  /* countbits.vhdl:86:31  */
  assign n32095_o = sum_r[64];
  /* countbits.vhdl:86:24  */
  assign n32097_o = {57'b000000000000000000000000000000000000000000000000000000000, n32095_o};
  /* countbits.vhdl:86:36  */
  assign n32098_o = {n32097_o, bitnum};
  /* countbits.vhdl:93:32  */
  assign n32102_o = pc8[31:28];
  /* countbits.vhdl:93:32  */
  assign n32103_o = pc8[27:24];
  /* countbits.vhdl:93:32  */
  assign n32104_o = pc8[23:20];
  /* countbits.vhdl:93:32  */
  assign n32105_o = pc8[19:16];
  /* countbits.vhdl:93:32  */
  assign n32106_o = pc8[15:12];
  /* countbits.vhdl:93:32  */
  assign n32107_o = pc8[11:8];
  /* countbits.vhdl:93:32  */
  assign n32108_o = pc8[7:4];
  /* countbits.vhdl:93:32  */
  assign n32109_o = pc8[3:0];
  assign n32112_o = {n32102_o, n32103_o, n32104_o, n32105_o, n32106_o, n32107_o, n32108_o, n32109_o};
  /* countbits.vhdl:103:40  */
  assign n32116_o = rs[0];
  /* countbits.vhdl:103:36  */
  assign n32118_o = {1'b0, n32116_o};
  /* countbits.vhdl:103:81  */
  assign n32119_o = rs[1];
  /* countbits.vhdl:103:77  */
  assign n32121_o = {1'b0, n32119_o};
  /* countbits.vhdl:103:62  */
  assign n32122_o = n32118_o + n32121_o;
  /* countbits.vhdl:103:40  */
  assign n32123_o = rs[2];
  /* countbits.vhdl:103:36  */
  assign n32125_o = {1'b0, n32123_o};
  /* countbits.vhdl:103:81  */
  assign n32126_o = rs[3];
  /* countbits.vhdl:103:77  */
  assign n32128_o = {1'b0, n32126_o};
  /* countbits.vhdl:103:62  */
  assign n32129_o = n32125_o + n32128_o;
  /* countbits.vhdl:103:40  */
  assign n32130_o = rs[4];
  /* countbits.vhdl:103:36  */
  assign n32132_o = {1'b0, n32130_o};
  /* countbits.vhdl:103:81  */
  assign n32133_o = rs[5];
  /* countbits.vhdl:103:77  */
  assign n32135_o = {1'b0, n32133_o};
  /* countbits.vhdl:103:62  */
  assign n32136_o = n32132_o + n32135_o;
  /* countbits.vhdl:103:40  */
  assign n32137_o = rs[6];
  /* countbits.vhdl:103:36  */
  assign n32139_o = {1'b0, n32137_o};
  /* countbits.vhdl:103:81  */
  assign n32140_o = rs[7];
  /* countbits.vhdl:103:77  */
  assign n32142_o = {1'b0, n32140_o};
  /* countbits.vhdl:103:62  */
  assign n32143_o = n32139_o + n32142_o;
  /* countbits.vhdl:103:40  */
  assign n32144_o = rs[8];
  /* countbits.vhdl:103:36  */
  assign n32146_o = {1'b0, n32144_o};
  /* countbits.vhdl:103:81  */
  assign n32147_o = rs[9];
  /* countbits.vhdl:103:77  */
  assign n32149_o = {1'b0, n32147_o};
  /* countbits.vhdl:103:62  */
  assign n32150_o = n32146_o + n32149_o;
  /* countbits.vhdl:103:40  */
  assign n32151_o = rs[10];
  /* countbits.vhdl:103:36  */
  assign n32153_o = {1'b0, n32151_o};
  /* countbits.vhdl:103:81  */
  assign n32154_o = rs[11];
  /* countbits.vhdl:103:77  */
  assign n32156_o = {1'b0, n32154_o};
  /* countbits.vhdl:103:62  */
  assign n32157_o = n32153_o + n32156_o;
  /* countbits.vhdl:103:40  */
  assign n32158_o = rs[12];
  /* countbits.vhdl:103:36  */
  assign n32160_o = {1'b0, n32158_o};
  /* countbits.vhdl:103:81  */
  assign n32161_o = rs[13];
  /* countbits.vhdl:103:77  */
  assign n32163_o = {1'b0, n32161_o};
  /* countbits.vhdl:103:62  */
  assign n32164_o = n32160_o + n32163_o;
  /* countbits.vhdl:103:40  */
  assign n32165_o = rs[14];
  /* countbits.vhdl:103:36  */
  assign n32167_o = {1'b0, n32165_o};
  /* countbits.vhdl:103:81  */
  assign n32168_o = rs[15];
  /* countbits.vhdl:103:77  */
  assign n32170_o = {1'b0, n32168_o};
  /* countbits.vhdl:103:62  */
  assign n32171_o = n32167_o + n32170_o;
  /* countbits.vhdl:103:40  */
  assign n32172_o = rs[16];
  /* countbits.vhdl:103:36  */
  assign n32174_o = {1'b0, n32172_o};
  /* countbits.vhdl:103:81  */
  assign n32175_o = rs[17];
  /* countbits.vhdl:103:77  */
  assign n32177_o = {1'b0, n32175_o};
  /* countbits.vhdl:103:62  */
  assign n32178_o = n32174_o + n32177_o;
  /* countbits.vhdl:103:40  */
  assign n32179_o = rs[18];
  /* countbits.vhdl:103:36  */
  assign n32181_o = {1'b0, n32179_o};
  /* countbits.vhdl:103:81  */
  assign n32182_o = rs[19];
  /* countbits.vhdl:103:77  */
  assign n32184_o = {1'b0, n32182_o};
  /* countbits.vhdl:103:62  */
  assign n32185_o = n32181_o + n32184_o;
  /* countbits.vhdl:103:40  */
  assign n32186_o = rs[20];
  /* countbits.vhdl:103:36  */
  assign n32188_o = {1'b0, n32186_o};
  /* countbits.vhdl:103:81  */
  assign n32189_o = rs[21];
  /* countbits.vhdl:103:77  */
  assign n32191_o = {1'b0, n32189_o};
  /* countbits.vhdl:103:62  */
  assign n32192_o = n32188_o + n32191_o;
  /* countbits.vhdl:103:40  */
  assign n32193_o = rs[22];
  /* countbits.vhdl:103:36  */
  assign n32195_o = {1'b0, n32193_o};
  /* countbits.vhdl:103:81  */
  assign n32196_o = rs[23];
  /* countbits.vhdl:103:77  */
  assign n32198_o = {1'b0, n32196_o};
  /* countbits.vhdl:103:62  */
  assign n32199_o = n32195_o + n32198_o;
  /* countbits.vhdl:103:40  */
  assign n32200_o = rs[24];
  /* countbits.vhdl:103:36  */
  assign n32202_o = {1'b0, n32200_o};
  /* countbits.vhdl:103:81  */
  assign n32203_o = rs[25];
  /* countbits.vhdl:103:77  */
  assign n32205_o = {1'b0, n32203_o};
  /* countbits.vhdl:103:62  */
  assign n32206_o = n32202_o + n32205_o;
  /* countbits.vhdl:103:40  */
  assign n32207_o = rs[26];
  /* countbits.vhdl:103:36  */
  assign n32209_o = {1'b0, n32207_o};
  /* countbits.vhdl:103:81  */
  assign n32210_o = rs[27];
  /* countbits.vhdl:103:77  */
  assign n32212_o = {1'b0, n32210_o};
  /* countbits.vhdl:103:62  */
  assign n32213_o = n32209_o + n32212_o;
  /* countbits.vhdl:103:40  */
  assign n32214_o = rs[28];
  /* countbits.vhdl:103:36  */
  assign n32216_o = {1'b0, n32214_o};
  /* countbits.vhdl:103:81  */
  assign n32217_o = rs[29];
  /* countbits.vhdl:103:77  */
  assign n32219_o = {1'b0, n32217_o};
  /* countbits.vhdl:103:62  */
  assign n32220_o = n32216_o + n32219_o;
  /* countbits.vhdl:103:40  */
  assign n32221_o = rs[30];
  /* countbits.vhdl:103:36  */
  assign n32223_o = {1'b0, n32221_o};
  /* countbits.vhdl:103:81  */
  assign n32224_o = rs[31];
  /* countbits.vhdl:103:77  */
  assign n32226_o = {1'b0, n32224_o};
  /* countbits.vhdl:103:62  */
  assign n32227_o = n32223_o + n32226_o;
  /* countbits.vhdl:103:40  */
  assign n32228_o = rs[32];
  /* countbits.vhdl:103:36  */
  assign n32230_o = {1'b0, n32228_o};
  /* countbits.vhdl:103:81  */
  assign n32231_o = rs[33];
  /* countbits.vhdl:103:77  */
  assign n32233_o = {1'b0, n32231_o};
  /* countbits.vhdl:103:62  */
  assign n32234_o = n32230_o + n32233_o;
  /* countbits.vhdl:103:40  */
  assign n32235_o = rs[34];
  /* countbits.vhdl:103:36  */
  assign n32237_o = {1'b0, n32235_o};
  /* countbits.vhdl:103:81  */
  assign n32238_o = rs[35];
  /* countbits.vhdl:103:77  */
  assign n32240_o = {1'b0, n32238_o};
  /* countbits.vhdl:103:62  */
  assign n32241_o = n32237_o + n32240_o;
  /* countbits.vhdl:103:40  */
  assign n32242_o = rs[36];
  /* countbits.vhdl:103:36  */
  assign n32244_o = {1'b0, n32242_o};
  /* countbits.vhdl:103:81  */
  assign n32245_o = rs[37];
  /* countbits.vhdl:103:77  */
  assign n32247_o = {1'b0, n32245_o};
  /* countbits.vhdl:103:62  */
  assign n32248_o = n32244_o + n32247_o;
  /* countbits.vhdl:103:40  */
  assign n32249_o = rs[38];
  /* countbits.vhdl:103:36  */
  assign n32251_o = {1'b0, n32249_o};
  /* countbits.vhdl:103:81  */
  assign n32252_o = rs[39];
  /* countbits.vhdl:103:77  */
  assign n32254_o = {1'b0, n32252_o};
  /* countbits.vhdl:103:62  */
  assign n32255_o = n32251_o + n32254_o;
  /* countbits.vhdl:103:40  */
  assign n32256_o = rs[40];
  /* countbits.vhdl:103:36  */
  assign n32258_o = {1'b0, n32256_o};
  /* countbits.vhdl:103:81  */
  assign n32259_o = rs[41];
  /* countbits.vhdl:103:77  */
  assign n32261_o = {1'b0, n32259_o};
  /* countbits.vhdl:103:62  */
  assign n32262_o = n32258_o + n32261_o;
  /* countbits.vhdl:103:40  */
  assign n32263_o = rs[42];
  /* countbits.vhdl:103:36  */
  assign n32265_o = {1'b0, n32263_o};
  /* countbits.vhdl:103:81  */
  assign n32266_o = rs[43];
  /* countbits.vhdl:103:77  */
  assign n32268_o = {1'b0, n32266_o};
  /* countbits.vhdl:103:62  */
  assign n32269_o = n32265_o + n32268_o;
  /* countbits.vhdl:103:40  */
  assign n32270_o = rs[44];
  /* countbits.vhdl:103:36  */
  assign n32272_o = {1'b0, n32270_o};
  /* countbits.vhdl:103:81  */
  assign n32273_o = rs[45];
  /* countbits.vhdl:103:77  */
  assign n32275_o = {1'b0, n32273_o};
  /* countbits.vhdl:103:62  */
  assign n32276_o = n32272_o + n32275_o;
  /* countbits.vhdl:103:40  */
  assign n32277_o = rs[46];
  /* countbits.vhdl:103:36  */
  assign n32279_o = {1'b0, n32277_o};
  /* countbits.vhdl:103:81  */
  assign n32280_o = rs[47];
  /* countbits.vhdl:103:77  */
  assign n32282_o = {1'b0, n32280_o};
  /* countbits.vhdl:103:62  */
  assign n32283_o = n32279_o + n32282_o;
  /* countbits.vhdl:103:40  */
  assign n32284_o = rs[48];
  /* countbits.vhdl:103:36  */
  assign n32286_o = {1'b0, n32284_o};
  /* countbits.vhdl:103:81  */
  assign n32287_o = rs[49];
  /* countbits.vhdl:103:77  */
  assign n32289_o = {1'b0, n32287_o};
  /* countbits.vhdl:103:62  */
  assign n32290_o = n32286_o + n32289_o;
  /* countbits.vhdl:103:40  */
  assign n32291_o = rs[50];
  /* countbits.vhdl:103:36  */
  assign n32293_o = {1'b0, n32291_o};
  /* countbits.vhdl:103:81  */
  assign n32294_o = rs[51];
  /* countbits.vhdl:103:77  */
  assign n32296_o = {1'b0, n32294_o};
  /* countbits.vhdl:103:62  */
  assign n32297_o = n32293_o + n32296_o;
  /* countbits.vhdl:103:40  */
  assign n32298_o = rs[52];
  /* countbits.vhdl:103:36  */
  assign n32300_o = {1'b0, n32298_o};
  /* countbits.vhdl:103:81  */
  assign n32301_o = rs[53];
  /* countbits.vhdl:103:77  */
  assign n32303_o = {1'b0, n32301_o};
  /* countbits.vhdl:103:62  */
  assign n32304_o = n32300_o + n32303_o;
  /* countbits.vhdl:103:40  */
  assign n32305_o = rs[54];
  /* countbits.vhdl:103:36  */
  assign n32307_o = {1'b0, n32305_o};
  /* countbits.vhdl:103:81  */
  assign n32308_o = rs[55];
  /* countbits.vhdl:103:77  */
  assign n32310_o = {1'b0, n32308_o};
  /* countbits.vhdl:103:62  */
  assign n32311_o = n32307_o + n32310_o;
  /* countbits.vhdl:103:40  */
  assign n32312_o = rs[56];
  /* countbits.vhdl:103:36  */
  assign n32314_o = {1'b0, n32312_o};
  /* countbits.vhdl:103:81  */
  assign n32315_o = rs[57];
  /* countbits.vhdl:103:77  */
  assign n32317_o = {1'b0, n32315_o};
  /* countbits.vhdl:103:62  */
  assign n32318_o = n32314_o + n32317_o;
  /* countbits.vhdl:103:40  */
  assign n32319_o = rs[58];
  /* countbits.vhdl:103:36  */
  assign n32321_o = {1'b0, n32319_o};
  /* countbits.vhdl:103:81  */
  assign n32322_o = rs[59];
  /* countbits.vhdl:103:77  */
  assign n32324_o = {1'b0, n32322_o};
  /* countbits.vhdl:103:62  */
  assign n32325_o = n32321_o + n32324_o;
  /* countbits.vhdl:103:40  */
  assign n32326_o = rs[60];
  /* countbits.vhdl:103:36  */
  assign n32328_o = {1'b0, n32326_o};
  /* countbits.vhdl:103:81  */
  assign n32329_o = rs[61];
  /* countbits.vhdl:103:77  */
  assign n32331_o = {1'b0, n32329_o};
  /* countbits.vhdl:103:62  */
  assign n32332_o = n32328_o + n32331_o;
  /* countbits.vhdl:103:40  */
  assign n32333_o = rs[62];
  /* countbits.vhdl:103:36  */
  assign n32335_o = {1'b0, n32333_o};
  /* countbits.vhdl:103:81  */
  assign n32336_o = rs[63];
  /* countbits.vhdl:103:77  */
  assign n32338_o = {1'b0, n32336_o};
  /* countbits.vhdl:103:62  */
  assign n32339_o = n32335_o + n32338_o;
  /* countbits.vhdl:106:33  */
  assign n32340_o = pc2[63:62];
  /* countbits.vhdl:106:28  */
  assign n32342_o = {1'b0, n32340_o};
  /* countbits.vhdl:106:54  */
  assign n32343_o = pc2[61:60];
  /* countbits.vhdl:106:49  */
  assign n32345_o = {1'b0, n32343_o};
  /* countbits.vhdl:106:42  */
  assign n32346_o = n32342_o + n32345_o;
  /* countbits.vhdl:106:33  */
  assign n32347_o = pc2[59:58];
  /* countbits.vhdl:106:28  */
  assign n32349_o = {1'b0, n32347_o};
  /* countbits.vhdl:106:54  */
  assign n32350_o = pc2[57:56];
  /* countbits.vhdl:106:49  */
  assign n32352_o = {1'b0, n32350_o};
  /* countbits.vhdl:106:42  */
  assign n32353_o = n32349_o + n32352_o;
  /* countbits.vhdl:106:33  */
  assign n32354_o = pc2[55:54];
  /* countbits.vhdl:106:28  */
  assign n32356_o = {1'b0, n32354_o};
  /* countbits.vhdl:106:54  */
  assign n32357_o = pc2[53:52];
  /* countbits.vhdl:106:49  */
  assign n32359_o = {1'b0, n32357_o};
  /* countbits.vhdl:106:42  */
  assign n32360_o = n32356_o + n32359_o;
  /* countbits.vhdl:106:33  */
  assign n32361_o = pc2[51:50];
  /* countbits.vhdl:106:28  */
  assign n32363_o = {1'b0, n32361_o};
  /* countbits.vhdl:106:54  */
  assign n32364_o = pc2[49:48];
  /* countbits.vhdl:106:49  */
  assign n32366_o = {1'b0, n32364_o};
  /* countbits.vhdl:106:42  */
  assign n32367_o = n32363_o + n32366_o;
  /* countbits.vhdl:106:33  */
  assign n32368_o = pc2[47:46];
  /* countbits.vhdl:106:28  */
  assign n32370_o = {1'b0, n32368_o};
  /* countbits.vhdl:106:54  */
  assign n32371_o = pc2[45:44];
  /* countbits.vhdl:106:49  */
  assign n32373_o = {1'b0, n32371_o};
  /* countbits.vhdl:106:42  */
  assign n32374_o = n32370_o + n32373_o;
  /* countbits.vhdl:106:33  */
  assign n32375_o = pc2[43:42];
  /* countbits.vhdl:106:28  */
  assign n32377_o = {1'b0, n32375_o};
  /* countbits.vhdl:106:54  */
  assign n32378_o = pc2[41:40];
  /* countbits.vhdl:106:49  */
  assign n32380_o = {1'b0, n32378_o};
  /* countbits.vhdl:106:42  */
  assign n32381_o = n32377_o + n32380_o;
  /* countbits.vhdl:106:33  */
  assign n32382_o = pc2[39:38];
  /* countbits.vhdl:106:28  */
  assign n32384_o = {1'b0, n32382_o};
  /* countbits.vhdl:106:54  */
  assign n32385_o = pc2[37:36];
  /* countbits.vhdl:106:49  */
  assign n32387_o = {1'b0, n32385_o};
  /* countbits.vhdl:106:42  */
  assign n32388_o = n32384_o + n32387_o;
  /* countbits.vhdl:106:33  */
  assign n32389_o = pc2[35:34];
  /* countbits.vhdl:106:28  */
  assign n32391_o = {1'b0, n32389_o};
  /* countbits.vhdl:106:54  */
  assign n32392_o = pc2[33:32];
  /* countbits.vhdl:106:49  */
  assign n32394_o = {1'b0, n32392_o};
  /* countbits.vhdl:106:42  */
  assign n32395_o = n32391_o + n32394_o;
  /* countbits.vhdl:106:33  */
  assign n32396_o = pc2[31:30];
  /* countbits.vhdl:106:28  */
  assign n32398_o = {1'b0, n32396_o};
  /* countbits.vhdl:106:54  */
  assign n32399_o = pc2[29:28];
  /* countbits.vhdl:106:49  */
  assign n32401_o = {1'b0, n32399_o};
  /* countbits.vhdl:106:42  */
  assign n32402_o = n32398_o + n32401_o;
  /* countbits.vhdl:106:33  */
  assign n32403_o = pc2[27:26];
  /* countbits.vhdl:106:28  */
  assign n32405_o = {1'b0, n32403_o};
  /* countbits.vhdl:106:54  */
  assign n32406_o = pc2[25:24];
  /* countbits.vhdl:106:49  */
  assign n32408_o = {1'b0, n32406_o};
  /* countbits.vhdl:106:42  */
  assign n32409_o = n32405_o + n32408_o;
  /* countbits.vhdl:106:33  */
  assign n32410_o = pc2[23:22];
  /* countbits.vhdl:106:28  */
  assign n32412_o = {1'b0, n32410_o};
  /* countbits.vhdl:106:54  */
  assign n32413_o = pc2[21:20];
  /* countbits.vhdl:106:49  */
  assign n32415_o = {1'b0, n32413_o};
  /* countbits.vhdl:106:42  */
  assign n32416_o = n32412_o + n32415_o;
  /* countbits.vhdl:106:33  */
  assign n32417_o = pc2[19:18];
  /* countbits.vhdl:106:28  */
  assign n32419_o = {1'b0, n32417_o};
  /* countbits.vhdl:106:54  */
  assign n32420_o = pc2[17:16];
  /* countbits.vhdl:106:49  */
  assign n32422_o = {1'b0, n32420_o};
  /* countbits.vhdl:106:42  */
  assign n32423_o = n32419_o + n32422_o;
  /* countbits.vhdl:106:33  */
  assign n32424_o = pc2[15:14];
  /* countbits.vhdl:106:28  */
  assign n32426_o = {1'b0, n32424_o};
  /* countbits.vhdl:106:54  */
  assign n32427_o = pc2[13:12];
  /* countbits.vhdl:106:49  */
  assign n32429_o = {1'b0, n32427_o};
  /* countbits.vhdl:106:42  */
  assign n32430_o = n32426_o + n32429_o;
  /* countbits.vhdl:106:33  */
  assign n32431_o = pc2[11:10];
  /* countbits.vhdl:106:28  */
  assign n32433_o = {1'b0, n32431_o};
  /* countbits.vhdl:106:54  */
  assign n32434_o = pc2[9:8];
  /* countbits.vhdl:106:49  */
  assign n32436_o = {1'b0, n32434_o};
  /* countbits.vhdl:106:42  */
  assign n32437_o = n32433_o + n32436_o;
  /* countbits.vhdl:106:33  */
  assign n32438_o = pc2[7:6];
  /* countbits.vhdl:106:28  */
  assign n32440_o = {1'b0, n32438_o};
  /* countbits.vhdl:106:54  */
  assign n32441_o = pc2[5:4];
  /* countbits.vhdl:106:49  */
  assign n32443_o = {1'b0, n32441_o};
  /* countbits.vhdl:106:42  */
  assign n32444_o = n32440_o + n32443_o;
  /* countbits.vhdl:106:33  */
  assign n32445_o = pc2[3:2];
  /* countbits.vhdl:106:28  */
  assign n32447_o = {1'b0, n32445_o};
  /* countbits.vhdl:106:54  */
  assign n32448_o = pc2[1:0];
  /* countbits.vhdl:106:49  */
  assign n32450_o = {1'b0, n32448_o};
  /* countbits.vhdl:106:42  */
  assign n32451_o = n32447_o + n32450_o;
  /* countbits.vhdl:109:33  */
  assign n32452_o = pc4[47:45];
  /* countbits.vhdl:109:28  */
  assign n32454_o = {1'b0, n32452_o};
  /* countbits.vhdl:109:54  */
  assign n32455_o = pc4[44:42];
  /* countbits.vhdl:109:49  */
  assign n32457_o = {1'b0, n32455_o};
  /* countbits.vhdl:109:42  */
  assign n32458_o = n32454_o + n32457_o;
  /* countbits.vhdl:109:33  */
  assign n32459_o = pc4[41:39];
  /* countbits.vhdl:109:28  */
  assign n32461_o = {1'b0, n32459_o};
  /* countbits.vhdl:109:54  */
  assign n32462_o = pc4[38:36];
  /* countbits.vhdl:109:49  */
  assign n32464_o = {1'b0, n32462_o};
  /* countbits.vhdl:109:42  */
  assign n32465_o = n32461_o + n32464_o;
  /* countbits.vhdl:109:33  */
  assign n32466_o = pc4[35:33];
  /* countbits.vhdl:109:28  */
  assign n32468_o = {1'b0, n32466_o};
  /* countbits.vhdl:109:54  */
  assign n32469_o = pc4[32:30];
  /* countbits.vhdl:109:49  */
  assign n32471_o = {1'b0, n32469_o};
  /* countbits.vhdl:109:42  */
  assign n32472_o = n32468_o + n32471_o;
  /* countbits.vhdl:109:33  */
  assign n32473_o = pc4[29:27];
  /* countbits.vhdl:109:28  */
  assign n32475_o = {1'b0, n32473_o};
  /* countbits.vhdl:109:54  */
  assign n32476_o = pc4[26:24];
  /* countbits.vhdl:109:49  */
  assign n32478_o = {1'b0, n32476_o};
  /* countbits.vhdl:109:42  */
  assign n32479_o = n32475_o + n32478_o;
  /* countbits.vhdl:109:33  */
  assign n32480_o = pc4[23:21];
  /* countbits.vhdl:109:28  */
  assign n32482_o = {1'b0, n32480_o};
  /* countbits.vhdl:109:54  */
  assign n32483_o = pc4[20:18];
  /* countbits.vhdl:109:49  */
  assign n32485_o = {1'b0, n32483_o};
  /* countbits.vhdl:109:42  */
  assign n32486_o = n32482_o + n32485_o;
  /* countbits.vhdl:109:33  */
  assign n32487_o = pc4[17:15];
  /* countbits.vhdl:109:28  */
  assign n32489_o = {1'b0, n32487_o};
  /* countbits.vhdl:109:54  */
  assign n32490_o = pc4[14:12];
  /* countbits.vhdl:109:49  */
  assign n32492_o = {1'b0, n32490_o};
  /* countbits.vhdl:109:42  */
  assign n32493_o = n32489_o + n32492_o;
  /* countbits.vhdl:109:33  */
  assign n32494_o = pc4[11:9];
  /* countbits.vhdl:109:28  */
  assign n32496_o = {1'b0, n32494_o};
  /* countbits.vhdl:109:54  */
  assign n32497_o = pc4[8:6];
  /* countbits.vhdl:109:49  */
  assign n32499_o = {1'b0, n32497_o};
  /* countbits.vhdl:109:42  */
  assign n32500_o = n32496_o + n32499_o;
  /* countbits.vhdl:109:33  */
  assign n32501_o = pc4[5:3];
  /* countbits.vhdl:109:28  */
  assign n32503_o = {1'b0, n32501_o};
  /* countbits.vhdl:109:54  */
  assign n32504_o = pc4[2:0];
  /* countbits.vhdl:109:49  */
  assign n32506_o = {1'b0, n32504_o};
  /* countbits.vhdl:109:42  */
  assign n32507_o = n32503_o + n32506_o;
  /* countbits.vhdl:114:37  */
  assign n32508_o = pc8_r[31:28];
  /* countbits.vhdl:114:30  */
  assign n32510_o = {2'b00, n32508_o};
  /* countbits.vhdl:114:61  */
  assign n32511_o = pc8_r[27:24];
  /* countbits.vhdl:114:54  */
  assign n32513_o = {2'b00, n32511_o};
  /* countbits.vhdl:114:46  */
  assign n32514_o = n32510_o + n32513_o;
  /* countbits.vhdl:115:37  */
  assign n32515_o = pc8_r[23:20];
  /* countbits.vhdl:115:30  */
  assign n32517_o = {2'b00, n32515_o};
  /* countbits.vhdl:114:74  */
  assign n32518_o = n32514_o + n32517_o;
  /* countbits.vhdl:115:65  */
  assign n32519_o = pc8_r[19:16];
  /* countbits.vhdl:115:58  */
  assign n32521_o = {2'b00, n32519_o};
  /* countbits.vhdl:115:50  */
  assign n32522_o = n32518_o + n32521_o;
  /* countbits.vhdl:114:37  */
  assign n32523_o = pc8_r[15:12];
  /* countbits.vhdl:114:30  */
  assign n32525_o = {2'b00, n32523_o};
  /* countbits.vhdl:114:61  */
  assign n32526_o = pc8_r[11:8];
  /* countbits.vhdl:114:54  */
  assign n32528_o = {2'b00, n32526_o};
  /* countbits.vhdl:114:46  */
  assign n32529_o = n32525_o + n32528_o;
  /* countbits.vhdl:115:37  */
  assign n32530_o = pc8_r[7:4];
  /* countbits.vhdl:115:30  */
  assign n32532_o = {2'b00, n32530_o};
  /* countbits.vhdl:114:74  */
  assign n32533_o = n32529_o + n32532_o;
  /* countbits.vhdl:115:65  */
  assign n32534_o = pc8_r[3:0];
  /* countbits.vhdl:115:58  */
  assign n32536_o = {2'b00, n32534_o};
  /* countbits.vhdl:115:50  */
  assign n32537_o = n32533_o + n32536_o;
  /* countbits.vhdl:119:18  */
  assign n32538_o = dlen_r[3:2];
  /* countbits.vhdl:119:31  */
  assign n32540_o = n32538_o == 2'b00;
  /* countbits.vhdl:122:74  */
  assign n32541_o = pc8_r[31:28];
  /* countbits.vhdl:122:74  */
  assign n32542_o = pc8_r[27:24];
  /* countbits.vhdl:122:74  */
  assign n32543_o = pc8_r[23:20];
  /* countbits.vhdl:122:74  */
  assign n32544_o = pc8_r[19:16];
  /* countbits.vhdl:122:74  */
  assign n32545_o = pc8_r[15:12];
  /* countbits.vhdl:122:74  */
  assign n32546_o = pc8_r[11:8];
  /* countbits.vhdl:122:74  */
  assign n32547_o = pc8_r[7:4];
  /* countbits.vhdl:122:74  */
  assign n32548_o = pc8_r[3:0];
  /* countbits.vhdl:124:21  */
  assign n32549_o = dlen_r[3];
  /* countbits.vhdl:124:25  */
  assign n32550_o = ~n32549_o;
  /* countbits.vhdl:127:75  */
  assign n32551_o = pc32[11:6];
  /* countbits.vhdl:127:75  */
  assign n32552_o = pc32[5:0];
  /* countbits.vhdl:130:64  */
  assign n32553_o = pc32[11:6];
  /* countbits.vhdl:130:58  */
  assign n32555_o = {1'b0, n32553_o};
  /* countbits.vhdl:130:82  */
  assign n32556_o = pc32[5:0];
  /* countbits.vhdl:130:76  */
  assign n32558_o = {1'b0, n32556_o};
  /* countbits.vhdl:130:69  */
  assign n32559_o = n32555_o + n32558_o;
  assign n32560_o = n32559_o[5:0];
  /* countbits.vhdl:124:9  */
  assign n32561_o = n32550_o ? n32551_o : n32560_o;
  assign n32562_o = n32559_o[6];
  /* countbits.vhdl:124:9  */
  assign n32564_o = n32550_o ? 1'b0 : n32562_o;
  /* countbits.vhdl:124:9  */
  assign n32566_o = n32550_o ? n32552_o : 6'b000000;
  assign n32567_o = {n32564_o, n32561_o};
  assign n32568_o = n32567_o[3:0];
  /* countbits.vhdl:119:9  */
  assign n32569_o = n32540_o ? n32541_o : n32568_o;
  assign n32570_o = n32567_o[6:4];
  /* countbits.vhdl:119:9  */
  assign n32572_o = n32540_o ? 3'b000 : n32570_o;
  /* countbits.vhdl:119:9  */
  assign n32574_o = n32540_o ? n32542_o : 4'b0000;
  /* countbits.vhdl:119:9  */
  assign n32576_o = n32540_o ? n32543_o : 4'b0000;
  /* countbits.vhdl:119:9  */
  assign n32578_o = n32540_o ? n32544_o : 4'b0000;
  assign n32579_o = n32566_o[3:0];
  /* countbits.vhdl:119:9  */
  assign n32580_o = n32540_o ? n32545_o : n32579_o;
  assign n32581_o = n32566_o[5:4];
  /* countbits.vhdl:119:9  */
  assign n32583_o = n32540_o ? 2'b00 : n32581_o;
  /* countbits.vhdl:119:9  */
  assign n32585_o = n32540_o ? n32546_o : 4'b0000;
  /* countbits.vhdl:119:9  */
  assign n32587_o = n32540_o ? n32547_o : 4'b0000;
  /* countbits.vhdl:119:9  */
  assign n32589_o = n32540_o ? n32548_o : 4'b0000;
  assign n32594_o = n32590_o[7];
  assign n32596_o = n32590_o[15:12];
  assign n32598_o = n32590_o[23:20];
  assign n32600_o = n32590_o[31:28];
  assign n32603_o = n32590_o[39:38];
  assign n32605_o = n32590_o[47:44];
  assign n32606_o = n32590_o[63:60];
  assign n32607_o = n32590_o[55:52];
  /* countbits.vhdl:134:32  */
  assign n32609_o = ~pcnt_r;
  /* countbits.vhdl:134:20  */
  assign n32610_o = n32609_o ? cntz : popcnt;
  /* countbits.vhdl:52:9  */
  always @(posedge clk)
    n32611_q <= inp;
  /* countbits.vhdl:52:9  */
  always @(posedge clk)
    n32612_q <= sum;
  /* countbits.vhdl:52:9  */
  assign n32613_o = {n32093_o, n32094_o};
  /* countbits.vhdl:91:9  */
  always @(posedge clk)
    n32614_q <= datalen;
  /* countbits.vhdl:91:9  */
  always @(posedge clk)
    n32615_q <= do_popcnt;
  /* countbits.vhdl:91:9  */
  assign n32616_o = {n32122_o, n32129_o, n32136_o, n32143_o, n32150_o, n32157_o, n32164_o, n32171_o, n32178_o, n32185_o, n32192_o, n32199_o, n32206_o, n32213_o, n32220_o, n32227_o, n32234_o, n32241_o, n32248_o, n32255_o, n32262_o, n32269_o, n32276_o, n32283_o, n32290_o, n32297_o, n32304_o, n32311_o, n32318_o, n32325_o, n32332_o, n32339_o};
  assign n32617_o = {n32346_o, n32353_o, n32360_o, n32367_o, n32374_o, n32381_o, n32388_o, n32395_o, n32402_o, n32409_o, n32416_o, n32423_o, n32430_o, n32437_o, n32444_o, n32451_o};
  assign n32618_o = {n32458_o, n32465_o, n32472_o, n32479_o, n32486_o, n32493_o, n32500_o, n32507_o};
  /* countbits.vhdl:91:9  */
  always @(posedge clk)
    n32619_q <= n32112_o;
  /* countbits.vhdl:91:9  */
  assign n32620_o = {n32522_o, n32537_o};
  assign n32621_o = {n32606_o, n32589_o, n32607_o, n32587_o, n32605_o, n32585_o, n32603_o, n32583_o, n32580_o, n32600_o, n32578_o, n32598_o, n32576_o, n32596_o, n32574_o, n32594_o, n32572_o, n32569_o};
endmodule

module logical
  (input  [63:0] rs,
   input  [63:0] rb,
   input  [5:0] op,
   input  invert_in,
   input  invert_out,
   input  [3:0] datalen,
   output [63:0] result);
  wire par0;
  wire par1;
  wire [63:0] parity;
  wire [7:0] permute;
  wire n28917_o;
  wire n28918_o;
  wire n28919_o;
  wire n28920_o;
  wire n28921_o;
  wire n28922_o;
  wire n28923_o;
  wire n28924_o;
  wire n28925_o;
  wire n28926_o;
  wire n28927_o;
  wire n28928_o;
  wire n28929_o;
  wire n28930_o;
  wire n28931_o;
  wire n28932_o;
  wire n28933_o;
  wire n28935_o;
  localparam [63:0] n28936_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire [30:0] n28938_o;
  wire [30:0] n28939_o;
  wire [1:0] n28940_o;
  wire n28942_o;
  wire [5:0] n28943_o;
  wire [5:0] n28944_o;
  wire n28949_o;
  wire [1:0] n28950_o;
  wire n28952_o;
  wire [5:0] n28953_o;
  wire [5:0] n28954_o;
  wire n28959_o;
  wire [1:0] n28960_o;
  wire n28962_o;
  wire [5:0] n28963_o;
  wire [5:0] n28964_o;
  wire n28969_o;
  wire [1:0] n28970_o;
  wire n28972_o;
  wire [5:0] n28973_o;
  wire [5:0] n28974_o;
  wire n28979_o;
  wire [1:0] n28980_o;
  wire n28982_o;
  wire [5:0] n28983_o;
  wire [5:0] n28984_o;
  wire n28989_o;
  wire [1:0] n28990_o;
  wire n28992_o;
  wire [5:0] n28993_o;
  wire [5:0] n28994_o;
  wire n28999_o;
  wire [1:0] n29000_o;
  wire n29002_o;
  wire [5:0] n29003_o;
  wire [5:0] n29004_o;
  wire n29009_o;
  wire [1:0] n29010_o;
  wire n29012_o;
  wire [5:0] n29013_o;
  wire [5:0] n29014_o;
  wire n29019_o;
  wire [63:0] n29020_o;
  wire [63:0] n29021_o;
  wire [63:0] n29022_o;
  wire n29024_o;
  wire [63:0] n29025_o;
  wire n29027_o;
  wire [63:0] n29028_o;
  wire [1:0] n29029_o;
  reg [63:0] n29030_o;
  wire [63:0] n29031_o;
  wire [63:0] n29032_o;
  wire n29034_o;
  wire n29036_o;
  wire n29037_o;
  wire n29039_o;
  wire n29040_o;
  wire n29042_o;
  wire [7:0] n29052_o;
  wire [7:0] n29053_o;
  wire n29059_o;
  wire [7:0] n29062_o;
  wire [7:0] n29067_o;
  wire [7:0] n29068_o;
  wire n29074_o;
  wire [7:0] n29077_o;
  wire [7:0] n29081_o;
  wire [7:0] n29082_o;
  wire n29088_o;
  wire [7:0] n29091_o;
  wire [7:0] n29095_o;
  wire [7:0] n29096_o;
  wire n29102_o;
  wire [7:0] n29105_o;
  wire [7:0] n29109_o;
  wire [7:0] n29110_o;
  wire n29116_o;
  wire [7:0] n29119_o;
  wire [7:0] n29123_o;
  wire [7:0] n29124_o;
  wire n29130_o;
  wire [7:0] n29133_o;
  wire [7:0] n29137_o;
  wire [7:0] n29138_o;
  wire n29144_o;
  wire [7:0] n29147_o;
  wire [7:0] n29151_o;
  wire [7:0] n29152_o;
  wire n29158_o;
  wire [7:0] n29161_o;
  wire [63:0] n29163_o;
  wire n29165_o;
  wire [63:0] n29166_o;
  wire n29168_o;
  wire n29169_o;
  wire [11:0] n29171_o;
  wire n29189_o;
  wire n29191_o;
  wire n29193_o;
  wire n29195_o;
  wire n29197_o;
  wire n29199_o;
  wire n29201_o;
  wire n29203_o;
  wire n29205_o;
  wire n29207_o;
  wire n29209_o;
  wire n29211_o;
  wire n29213_o;
  wire n29214_o;
  wire n29215_o;
  wire n29216_o;
  wire n29217_o;
  wire n29218_o;
  wire n29219_o;
  wire n29220_o;
  wire n29221_o;
  wire n29222_o;
  wire n29223_o;
  wire n29226_o;
  wire n29227_o;
  wire n29228_o;
  wire n29229_o;
  wire n29230_o;
  wire n29231_o;
  wire n29232_o;
  wire n29233_o;
  wire n29234_o;
  wire n29235_o;
  wire n29236_o;
  wire n29239_o;
  wire n29240_o;
  wire n29241_o;
  wire n29242_o;
  wire n29243_o;
  wire n29244_o;
  wire n29245_o;
  wire n29246_o;
  wire n29247_o;
  wire n29248_o;
  wire n29249_o;
  wire n29250_o;
  wire n29251_o;
  wire n29252_o;
  wire n29253_o;
  wire n29254_o;
  wire n29255_o;
  wire n29257_o;
  wire n29258_o;
  wire n29259_o;
  wire n29260_o;
  wire n29261_o;
  wire n29262_o;
  wire n29263_o;
  wire n29264_o;
  wire n29265_o;
  wire n29266_o;
  wire n29267_o;
  wire n29268_o;
  wire n29269_o;
  wire n29270_o;
  wire n29271_o;
  wire n29272_o;
  wire n29273_o;
  wire n29276_o;
  wire n29277_o;
  wire n29279_o;
  wire n29280_o;
  wire n29281_o;
  wire n29282_o;
  wire n29283_o;
  wire n29284_o;
  wire n29285_o;
  wire n29287_o;
  wire n29288_o;
  wire n29289_o;
  wire n29290_o;
  wire n29291_o;
  wire n29292_o;
  wire n29293_o;
  wire [9:0] n29295_o;
  wire [21:0] n29297_o;
  wire [11:0] n29299_o;
  wire n29317_o;
  wire n29319_o;
  wire n29321_o;
  wire n29323_o;
  wire n29325_o;
  wire n29327_o;
  wire n29329_o;
  wire n29331_o;
  wire n29333_o;
  wire n29335_o;
  wire n29337_o;
  wire n29339_o;
  wire n29341_o;
  wire n29342_o;
  wire n29343_o;
  wire n29344_o;
  wire n29345_o;
  wire n29346_o;
  wire n29347_o;
  wire n29348_o;
  wire n29349_o;
  wire n29350_o;
  wire n29351_o;
  wire n29354_o;
  wire n29355_o;
  wire n29356_o;
  wire n29357_o;
  wire n29358_o;
  wire n29359_o;
  wire n29360_o;
  wire n29361_o;
  wire n29362_o;
  wire n29363_o;
  wire n29364_o;
  wire n29367_o;
  wire n29368_o;
  wire n29369_o;
  wire n29370_o;
  wire n29371_o;
  wire n29372_o;
  wire n29373_o;
  wire n29374_o;
  wire n29375_o;
  wire n29376_o;
  wire n29377_o;
  wire n29378_o;
  wire n29379_o;
  wire n29380_o;
  wire n29381_o;
  wire n29382_o;
  wire n29383_o;
  wire n29385_o;
  wire n29386_o;
  wire n29387_o;
  wire n29388_o;
  wire n29389_o;
  wire n29390_o;
  wire n29391_o;
  wire n29392_o;
  wire n29393_o;
  wire n29394_o;
  wire n29395_o;
  wire n29396_o;
  wire n29397_o;
  wire n29398_o;
  wire n29399_o;
  wire n29400_o;
  wire n29401_o;
  wire n29404_o;
  wire n29405_o;
  wire n29407_o;
  wire n29408_o;
  wire n29409_o;
  wire n29410_o;
  wire n29411_o;
  wire n29412_o;
  wire n29413_o;
  wire n29415_o;
  wire n29416_o;
  wire n29417_o;
  wire n29418_o;
  wire n29419_o;
  wire n29420_o;
  wire n29421_o;
  wire [9:0] n29423_o;
  wire [31:0] n29424_o;
  wire [43:0] n29426_o;
  wire [11:0] n29428_o;
  wire n29446_o;
  wire n29448_o;
  wire n29450_o;
  wire n29452_o;
  wire n29454_o;
  wire n29456_o;
  wire n29458_o;
  wire n29460_o;
  wire n29462_o;
  wire n29464_o;
  wire n29466_o;
  wire n29468_o;
  wire n29470_o;
  wire n29471_o;
  wire n29472_o;
  wire n29473_o;
  wire n29474_o;
  wire n29475_o;
  wire n29476_o;
  wire n29477_o;
  wire n29478_o;
  wire n29479_o;
  wire n29480_o;
  wire n29483_o;
  wire n29484_o;
  wire n29485_o;
  wire n29486_o;
  wire n29487_o;
  wire n29488_o;
  wire n29489_o;
  wire n29490_o;
  wire n29491_o;
  wire n29492_o;
  wire n29493_o;
  wire n29496_o;
  wire n29497_o;
  wire n29498_o;
  wire n29499_o;
  wire n29500_o;
  wire n29501_o;
  wire n29502_o;
  wire n29503_o;
  wire n29504_o;
  wire n29505_o;
  wire n29506_o;
  wire n29507_o;
  wire n29508_o;
  wire n29509_o;
  wire n29510_o;
  wire n29511_o;
  wire n29512_o;
  wire n29514_o;
  wire n29515_o;
  wire n29516_o;
  wire n29517_o;
  wire n29518_o;
  wire n29519_o;
  wire n29520_o;
  wire n29521_o;
  wire n29522_o;
  wire n29523_o;
  wire n29524_o;
  wire n29525_o;
  wire n29526_o;
  wire n29527_o;
  wire n29528_o;
  wire n29529_o;
  wire n29530_o;
  wire n29533_o;
  wire n29534_o;
  wire n29536_o;
  wire n29537_o;
  wire n29538_o;
  wire n29539_o;
  wire n29540_o;
  wire n29541_o;
  wire n29542_o;
  wire n29544_o;
  wire n29545_o;
  wire n29546_o;
  wire n29547_o;
  wire n29548_o;
  wire n29549_o;
  wire n29550_o;
  wire [9:0] n29552_o;
  wire [53:0] n29553_o;
  wire [11:0] n29555_o;
  wire n29573_o;
  wire n29575_o;
  wire n29577_o;
  wire n29579_o;
  wire n29581_o;
  wire n29583_o;
  wire n29585_o;
  wire n29587_o;
  wire n29589_o;
  wire n29591_o;
  wire n29593_o;
  wire n29595_o;
  wire n29597_o;
  wire n29598_o;
  wire n29599_o;
  wire n29600_o;
  wire n29601_o;
  wire n29602_o;
  wire n29603_o;
  wire n29604_o;
  wire n29605_o;
  wire n29606_o;
  wire n29607_o;
  wire n29610_o;
  wire n29611_o;
  wire n29612_o;
  wire n29613_o;
  wire n29614_o;
  wire n29615_o;
  wire n29616_o;
  wire n29617_o;
  wire n29618_o;
  wire n29619_o;
  wire n29620_o;
  wire n29623_o;
  wire n29624_o;
  wire n29625_o;
  wire n29626_o;
  wire n29627_o;
  wire n29628_o;
  wire n29629_o;
  wire n29630_o;
  wire n29631_o;
  wire n29632_o;
  wire n29633_o;
  wire n29634_o;
  wire n29635_o;
  wire n29636_o;
  wire n29637_o;
  wire n29638_o;
  wire n29639_o;
  wire n29641_o;
  wire n29642_o;
  wire n29643_o;
  wire n29644_o;
  wire n29645_o;
  wire n29646_o;
  wire n29647_o;
  wire n29648_o;
  wire n29649_o;
  wire n29650_o;
  wire n29651_o;
  wire n29652_o;
  wire n29653_o;
  wire n29654_o;
  wire n29655_o;
  wire n29656_o;
  wire n29657_o;
  wire n29660_o;
  wire n29661_o;
  wire n29663_o;
  wire n29664_o;
  wire n29665_o;
  wire n29666_o;
  wire n29667_o;
  wire n29668_o;
  wire n29669_o;
  wire n29671_o;
  wire n29672_o;
  wire n29673_o;
  wire n29674_o;
  wire n29675_o;
  wire n29676_o;
  wire n29677_o;
  wire [9:0] n29679_o;
  wire [63:0] n29680_o;
  wire [9:0] n29682_o;
  wire n29698_o;
  wire n29700_o;
  wire n29702_o;
  wire n29704_o;
  wire n29706_o;
  wire n29708_o;
  wire n29710_o;
  wire n29712_o;
  wire n29714_o;
  wire n29716_o;
  wire n29718_o;
  wire n29719_o;
  wire n29720_o;
  wire n29721_o;
  wire n29722_o;
  wire n29723_o;
  wire n29724_o;
  wire n29725_o;
  wire n29726_o;
  wire n29727_o;
  wire n29728_o;
  wire n29731_o;
  wire n29732_o;
  wire n29733_o;
  wire n29734_o;
  wire n29735_o;
  wire n29736_o;
  wire n29737_o;
  wire n29738_o;
  wire n29739_o;
  wire n29740_o;
  wire n29742_o;
  wire n29743_o;
  wire n29744_o;
  wire n29745_o;
  wire n29746_o;
  wire n29747_o;
  wire n29748_o;
  wire n29749_o;
  wire n29750_o;
  wire n29751_o;
  wire n29754_o;
  wire n29755_o;
  wire n29756_o;
  wire n29757_o;
  wire n29758_o;
  wire n29759_o;
  wire n29760_o;
  wire n29761_o;
  wire n29762_o;
  wire n29763_o;
  wire n29764_o;
  wire n29765_o;
  wire n29767_o;
  wire n29768_o;
  wire n29769_o;
  wire n29770_o;
  wire n29771_o;
  wire n29772_o;
  wire n29773_o;
  wire n29774_o;
  wire n29775_o;
  wire n29776_o;
  wire n29777_o;
  wire n29778_o;
  wire n29779_o;
  wire n29781_o;
  wire n29782_o;
  wire n29783_o;
  wire n29784_o;
  wire n29785_o;
  wire n29786_o;
  wire n29787_o;
  wire n29788_o;
  wire n29789_o;
  wire n29790_o;
  wire n29791_o;
  wire n29792_o;
  wire n29793_o;
  wire n29796_o;
  wire n29797_o;
  wire n29798_o;
  wire n29799_o;
  wire n29800_o;
  wire n29801_o;
  wire n29802_o;
  wire n29803_o;
  wire n29804_o;
  wire n29805_o;
  wire n29806_o;
  wire n29807_o;
  wire n29809_o;
  wire n29810_o;
  wire n29811_o;
  wire n29812_o;
  wire n29813_o;
  wire n29814_o;
  wire n29815_o;
  wire n29816_o;
  wire n29817_o;
  wire n29818_o;
  wire n29819_o;
  wire n29820_o;
  wire n29821_o;
  wire n29822_o;
  wire n29823_o;
  wire n29824_o;
  wire n29825_o;
  wire n29826_o;
  wire n29827_o;
  wire n29829_o;
  wire n29830_o;
  wire n29831_o;
  wire n29832_o;
  wire n29833_o;
  wire n29834_o;
  wire n29835_o;
  wire n29836_o;
  wire n29837_o;
  wire n29838_o;
  wire n29839_o;
  wire n29840_o;
  wire n29841_o;
  wire n29842_o;
  wire n29843_o;
  wire n29844_o;
  wire n29845_o;
  wire n29846_o;
  wire n29847_o;
  wire [11:0] n29849_o;
  wire [19:0] n29851_o;
  wire [9:0] n29853_o;
  wire n29869_o;
  wire n29871_o;
  wire n29873_o;
  wire n29875_o;
  wire n29877_o;
  wire n29879_o;
  wire n29881_o;
  wire n29883_o;
  wire n29885_o;
  wire n29887_o;
  wire n29889_o;
  wire n29890_o;
  wire n29891_o;
  wire n29892_o;
  wire n29893_o;
  wire n29894_o;
  wire n29895_o;
  wire n29896_o;
  wire n29897_o;
  wire n29898_o;
  wire n29899_o;
  wire n29902_o;
  wire n29903_o;
  wire n29904_o;
  wire n29905_o;
  wire n29906_o;
  wire n29907_o;
  wire n29908_o;
  wire n29909_o;
  wire n29910_o;
  wire n29911_o;
  wire n29913_o;
  wire n29914_o;
  wire n29915_o;
  wire n29916_o;
  wire n29917_o;
  wire n29918_o;
  wire n29919_o;
  wire n29920_o;
  wire n29921_o;
  wire n29922_o;
  wire n29925_o;
  wire n29926_o;
  wire n29927_o;
  wire n29928_o;
  wire n29929_o;
  wire n29930_o;
  wire n29931_o;
  wire n29932_o;
  wire n29933_o;
  wire n29934_o;
  wire n29935_o;
  wire n29936_o;
  wire n29938_o;
  wire n29939_o;
  wire n29940_o;
  wire n29941_o;
  wire n29942_o;
  wire n29943_o;
  wire n29944_o;
  wire n29945_o;
  wire n29946_o;
  wire n29947_o;
  wire n29948_o;
  wire n29949_o;
  wire n29950_o;
  wire n29952_o;
  wire n29953_o;
  wire n29954_o;
  wire n29955_o;
  wire n29956_o;
  wire n29957_o;
  wire n29958_o;
  wire n29959_o;
  wire n29960_o;
  wire n29961_o;
  wire n29962_o;
  wire n29963_o;
  wire n29964_o;
  wire n29967_o;
  wire n29968_o;
  wire n29969_o;
  wire n29970_o;
  wire n29971_o;
  wire n29972_o;
  wire n29973_o;
  wire n29974_o;
  wire n29975_o;
  wire n29976_o;
  wire n29977_o;
  wire n29978_o;
  wire n29980_o;
  wire n29981_o;
  wire n29982_o;
  wire n29983_o;
  wire n29984_o;
  wire n29985_o;
  wire n29986_o;
  wire n29987_o;
  wire n29988_o;
  wire n29989_o;
  wire n29990_o;
  wire n29991_o;
  wire n29992_o;
  wire n29993_o;
  wire n29994_o;
  wire n29995_o;
  wire n29996_o;
  wire n29997_o;
  wire n29998_o;
  wire n30000_o;
  wire n30001_o;
  wire n30002_o;
  wire n30003_o;
  wire n30004_o;
  wire n30005_o;
  wire n30006_o;
  wire n30007_o;
  wire n30008_o;
  wire n30009_o;
  wire n30010_o;
  wire n30011_o;
  wire n30012_o;
  wire n30013_o;
  wire n30014_o;
  wire n30015_o;
  wire n30016_o;
  wire n30017_o;
  wire n30018_o;
  wire [11:0] n30020_o;
  wire [31:0] n30021_o;
  wire [39:0] n30023_o;
  wire [9:0] n30025_o;
  wire n30041_o;
  wire n30043_o;
  wire n30045_o;
  wire n30047_o;
  wire n30049_o;
  wire n30051_o;
  wire n30053_o;
  wire n30055_o;
  wire n30057_o;
  wire n30059_o;
  wire n30061_o;
  wire n30062_o;
  wire n30063_o;
  wire n30064_o;
  wire n30065_o;
  wire n30066_o;
  wire n30067_o;
  wire n30068_o;
  wire n30069_o;
  wire n30070_o;
  wire n30071_o;
  wire n30074_o;
  wire n30075_o;
  wire n30076_o;
  wire n30077_o;
  wire n30078_o;
  wire n30079_o;
  wire n30080_o;
  wire n30081_o;
  wire n30082_o;
  wire n30083_o;
  wire n30085_o;
  wire n30086_o;
  wire n30087_o;
  wire n30088_o;
  wire n30089_o;
  wire n30090_o;
  wire n30091_o;
  wire n30092_o;
  wire n30093_o;
  wire n30094_o;
  wire n30097_o;
  wire n30098_o;
  wire n30099_o;
  wire n30100_o;
  wire n30101_o;
  wire n30102_o;
  wire n30103_o;
  wire n30104_o;
  wire n30105_o;
  wire n30106_o;
  wire n30107_o;
  wire n30108_o;
  wire n30110_o;
  wire n30111_o;
  wire n30112_o;
  wire n30113_o;
  wire n30114_o;
  wire n30115_o;
  wire n30116_o;
  wire n30117_o;
  wire n30118_o;
  wire n30119_o;
  wire n30120_o;
  wire n30121_o;
  wire n30122_o;
  wire n30124_o;
  wire n30125_o;
  wire n30126_o;
  wire n30127_o;
  wire n30128_o;
  wire n30129_o;
  wire n30130_o;
  wire n30131_o;
  wire n30132_o;
  wire n30133_o;
  wire n30134_o;
  wire n30135_o;
  wire n30136_o;
  wire n30139_o;
  wire n30140_o;
  wire n30141_o;
  wire n30142_o;
  wire n30143_o;
  wire n30144_o;
  wire n30145_o;
  wire n30146_o;
  wire n30147_o;
  wire n30148_o;
  wire n30149_o;
  wire n30150_o;
  wire n30152_o;
  wire n30153_o;
  wire n30154_o;
  wire n30155_o;
  wire n30156_o;
  wire n30157_o;
  wire n30158_o;
  wire n30159_o;
  wire n30160_o;
  wire n30161_o;
  wire n30162_o;
  wire n30163_o;
  wire n30164_o;
  wire n30165_o;
  wire n30166_o;
  wire n30167_o;
  wire n30168_o;
  wire n30169_o;
  wire n30170_o;
  wire n30172_o;
  wire n30173_o;
  wire n30174_o;
  wire n30175_o;
  wire n30176_o;
  wire n30177_o;
  wire n30178_o;
  wire n30179_o;
  wire n30180_o;
  wire n30181_o;
  wire n30182_o;
  wire n30183_o;
  wire n30184_o;
  wire n30185_o;
  wire n30186_o;
  wire n30187_o;
  wire n30188_o;
  wire n30189_o;
  wire n30190_o;
  wire [11:0] n30192_o;
  wire [51:0] n30193_o;
  wire [9:0] n30195_o;
  wire n30211_o;
  wire n30213_o;
  wire n30215_o;
  wire n30217_o;
  wire n30219_o;
  wire n30221_o;
  wire n30223_o;
  wire n30225_o;
  wire n30227_o;
  wire n30229_o;
  wire n30231_o;
  wire n30232_o;
  wire n30233_o;
  wire n30234_o;
  wire n30235_o;
  wire n30236_o;
  wire n30237_o;
  wire n30238_o;
  wire n30239_o;
  wire n30240_o;
  wire n30241_o;
  wire n30244_o;
  wire n30245_o;
  wire n30246_o;
  wire n30247_o;
  wire n30248_o;
  wire n30249_o;
  wire n30250_o;
  wire n30251_o;
  wire n30252_o;
  wire n30253_o;
  wire n30255_o;
  wire n30256_o;
  wire n30257_o;
  wire n30258_o;
  wire n30259_o;
  wire n30260_o;
  wire n30261_o;
  wire n30262_o;
  wire n30263_o;
  wire n30264_o;
  wire n30267_o;
  wire n30268_o;
  wire n30269_o;
  wire n30270_o;
  wire n30271_o;
  wire n30272_o;
  wire n30273_o;
  wire n30274_o;
  wire n30275_o;
  wire n30276_o;
  wire n30277_o;
  wire n30278_o;
  wire n30280_o;
  wire n30281_o;
  wire n30282_o;
  wire n30283_o;
  wire n30284_o;
  wire n30285_o;
  wire n30286_o;
  wire n30287_o;
  wire n30288_o;
  wire n30289_o;
  wire n30290_o;
  wire n30291_o;
  wire n30292_o;
  wire n30294_o;
  wire n30295_o;
  wire n30296_o;
  wire n30297_o;
  wire n30298_o;
  wire n30299_o;
  wire n30300_o;
  wire n30301_o;
  wire n30302_o;
  wire n30303_o;
  wire n30304_o;
  wire n30305_o;
  wire n30306_o;
  wire n30309_o;
  wire n30310_o;
  wire n30311_o;
  wire n30312_o;
  wire n30313_o;
  wire n30314_o;
  wire n30315_o;
  wire n30316_o;
  wire n30317_o;
  wire n30318_o;
  wire n30319_o;
  wire n30320_o;
  wire n30322_o;
  wire n30323_o;
  wire n30324_o;
  wire n30325_o;
  wire n30326_o;
  wire n30327_o;
  wire n30328_o;
  wire n30329_o;
  wire n30330_o;
  wire n30331_o;
  wire n30332_o;
  wire n30333_o;
  wire n30334_o;
  wire n30335_o;
  wire n30336_o;
  wire n30337_o;
  wire n30338_o;
  wire n30339_o;
  wire n30340_o;
  wire n30342_o;
  wire n30343_o;
  wire n30344_o;
  wire n30345_o;
  wire n30346_o;
  wire n30347_o;
  wire n30348_o;
  wire n30349_o;
  wire n30350_o;
  wire n30351_o;
  wire n30352_o;
  wire n30353_o;
  wire n30354_o;
  wire n30355_o;
  wire n30356_o;
  wire n30357_o;
  wire n30358_o;
  wire n30359_o;
  wire n30360_o;
  wire [11:0] n30362_o;
  wire [63:0] n30363_o;
  wire [63:0] n30364_o;
  wire n30366_o;
  wire n30367_o;
  wire n30368_o;
  wire n30369_o;
  wire n30370_o;
  wire n30371_o;
  wire n30372_o;
  wire n30373_o;
  wire n30374_o;
  wire n30375_o;
  wire n30376_o;
  wire n30377_o;
  wire [3:0] n30378_o;
  wire [3:0] n30379_o;
  wire [3:0] n30380_o;
  wire [3:0] n30381_o;
  wire [3:0] n30382_o;
  wire [3:0] n30383_o;
  wire [3:0] n30384_o;
  wire [3:0] n30385_o;
  wire [3:0] n30386_o;
  wire [3:0] n30387_o;
  wire [3:0] n30388_o;
  wire [3:0] n30389_o;
  wire [3:0] n30390_o;
  wire [3:0] n30391_o;
  wire [3:0] n30392_o;
  wire [3:0] n30393_o;
  wire [15:0] n30394_o;
  wire [15:0] n30395_o;
  wire [15:0] n30396_o;
  wire [15:0] n30397_o;
  wire [63:0] n30398_o;
  wire n30399_o;
  wire [15:0] n30400_o;
  wire [15:0] n30401_o;
  wire [15:0] n30402_o;
  wire [31:0] n30403_o;
  wire n30405_o;
  wire n30406_o;
  wire n30407_o;
  wire [7:0] n30408_o;
  wire [7:0] n30409_o;
  wire [7:0] n30410_o;
  wire [7:0] n30412_o;
  wire n30414_o;
  wire [5:0] n30415_o;
  wire [7:0] n30416_o;
  wire [7:0] n30417_o;
  wire [7:0] n30418_o;
  wire [7:0] n30419_o;
  wire [7:0] n30420_o;
  wire [7:0] n30421_o;
  reg [7:0] n30422_o;
  wire [7:0] n30423_o;
  wire [7:0] n30424_o;
  wire [7:0] n30425_o;
  wire [7:0] n30426_o;
  wire [7:0] n30427_o;
  wire [7:0] n30428_o;
  reg [7:0] n30429_o;
  wire [15:0] n30430_o;
  wire [15:0] n30431_o;
  wire [15:0] n30432_o;
  wire [15:0] n30433_o;
  wire [15:0] n30434_o;
  wire [15:0] n30435_o;
  reg [15:0] n30436_o;
  wire [31:0] n30437_o;
  wire [31:0] n30438_o;
  wire [31:0] n30439_o;
  wire [31:0] n30440_o;
  wire [31:0] n30441_o;
  wire [31:0] n30442_o;
  reg [31:0] n30443_o;
  wire [63:0] n30445_o;
  wire [63:0] n30449_o;
  wire [7:0] n30450_o;
  wire n30451_o;
  wire n30452_o;
  wire n30453_o;
  wire n30454_o;
  wire n30455_o;
  wire n30456_o;
  wire n30457_o;
  wire n30458_o;
  wire n30459_o;
  wire n30460_o;
  wire n30461_o;
  wire n30462_o;
  wire n30463_o;
  wire n30464_o;
  wire n30465_o;
  wire n30466_o;
  wire n30467_o;
  wire n30468_o;
  wire n30469_o;
  wire n30470_o;
  wire n30471_o;
  wire n30472_o;
  wire n30473_o;
  wire n30474_o;
  wire n30475_o;
  wire n30476_o;
  wire n30477_o;
  wire n30478_o;
  wire n30479_o;
  wire n30480_o;
  wire n30481_o;
  wire n30482_o;
  wire n30483_o;
  wire n30484_o;
  wire n30485_o;
  wire n30486_o;
  wire n30487_o;
  wire n30488_o;
  wire n30489_o;
  wire n30490_o;
  wire n30491_o;
  wire n30492_o;
  wire n30493_o;
  wire n30494_o;
  wire n30495_o;
  wire n30496_o;
  wire n30497_o;
  wire n30498_o;
  wire n30499_o;
  wire n30500_o;
  wire n30501_o;
  wire n30502_o;
  wire n30503_o;
  wire n30504_o;
  wire n30505_o;
  wire n30506_o;
  wire n30507_o;
  wire n30508_o;
  wire n30509_o;
  wire n30510_o;
  wire n30511_o;
  wire n30512_o;
  wire n30513_o;
  wire n30514_o;
  wire [1:0] n30515_o;
  reg n30516_o;
  wire [1:0] n30517_o;
  reg n30518_o;
  wire [1:0] n30519_o;
  reg n30520_o;
  wire [1:0] n30521_o;
  reg n30522_o;
  wire [1:0] n30523_o;
  reg n30524_o;
  wire [1:0] n30525_o;
  reg n30526_o;
  wire [1:0] n30527_o;
  reg n30528_o;
  wire [1:0] n30529_o;
  reg n30530_o;
  wire [1:0] n30531_o;
  reg n30532_o;
  wire [1:0] n30533_o;
  reg n30534_o;
  wire [1:0] n30535_o;
  reg n30536_o;
  wire [1:0] n30537_o;
  reg n30538_o;
  wire [1:0] n30539_o;
  reg n30540_o;
  wire [1:0] n30541_o;
  reg n30542_o;
  wire [1:0] n30543_o;
  reg n30544_o;
  wire [1:0] n30545_o;
  reg n30546_o;
  wire [1:0] n30547_o;
  reg n30548_o;
  wire [1:0] n30549_o;
  reg n30550_o;
  wire [1:0] n30551_o;
  reg n30552_o;
  wire [1:0] n30553_o;
  reg n30554_o;
  wire [1:0] n30555_o;
  reg n30556_o;
  wire n30557_o;
  wire n30558_o;
  wire n30559_o;
  wire n30560_o;
  wire n30561_o;
  wire n30562_o;
  wire n30563_o;
  wire n30564_o;
  wire n30565_o;
  wire n30566_o;
  wire n30567_o;
  wire n30568_o;
  wire n30569_o;
  wire n30570_o;
  wire n30571_o;
  wire n30572_o;
  wire n30573_o;
  wire n30574_o;
  wire n30575_o;
  wire n30576_o;
  wire n30577_o;
  wire n30578_o;
  wire n30579_o;
  wire n30580_o;
  wire n30581_o;
  wire n30582_o;
  wire n30583_o;
  wire n30584_o;
  wire n30585_o;
  wire n30586_o;
  wire n30587_o;
  wire n30588_o;
  wire n30589_o;
  wire n30590_o;
  wire n30591_o;
  wire n30592_o;
  wire n30593_o;
  wire n30594_o;
  wire n30595_o;
  wire n30596_o;
  wire n30597_o;
  wire n30598_o;
  wire n30599_o;
  wire n30600_o;
  wire n30601_o;
  wire n30602_o;
  wire n30603_o;
  wire n30604_o;
  wire n30605_o;
  wire n30606_o;
  wire n30607_o;
  wire n30608_o;
  wire n30609_o;
  wire n30610_o;
  wire n30611_o;
  wire n30612_o;
  wire n30613_o;
  wire n30614_o;
  wire n30615_o;
  wire n30616_o;
  wire n30617_o;
  wire n30618_o;
  wire n30619_o;
  wire n30620_o;
  wire [1:0] n30621_o;
  reg n30622_o;
  wire [1:0] n30623_o;
  reg n30624_o;
  wire [1:0] n30625_o;
  reg n30626_o;
  wire [1:0] n30627_o;
  reg n30628_o;
  wire [1:0] n30629_o;
  reg n30630_o;
  wire [1:0] n30631_o;
  reg n30632_o;
  wire [1:0] n30633_o;
  reg n30634_o;
  wire [1:0] n30635_o;
  reg n30636_o;
  wire [1:0] n30637_o;
  reg n30638_o;
  wire [1:0] n30639_o;
  reg n30640_o;
  wire [1:0] n30641_o;
  reg n30642_o;
  wire [1:0] n30643_o;
  reg n30644_o;
  wire [1:0] n30645_o;
  reg n30646_o;
  wire [1:0] n30647_o;
  reg n30648_o;
  wire [1:0] n30649_o;
  reg n30650_o;
  wire [1:0] n30651_o;
  reg n30652_o;
  wire [1:0] n30653_o;
  reg n30654_o;
  wire [1:0] n30655_o;
  reg n30656_o;
  wire [1:0] n30657_o;
  reg n30658_o;
  wire [1:0] n30659_o;
  reg n30660_o;
  wire [1:0] n30661_o;
  reg n30662_o;
  wire n30663_o;
  wire n30664_o;
  wire n30665_o;
  wire n30666_o;
  wire n30667_o;
  wire n30668_o;
  wire n30669_o;
  wire n30670_o;
  wire n30671_o;
  wire n30672_o;
  wire n30673_o;
  wire n30674_o;
  wire n30675_o;
  wire n30676_o;
  wire n30677_o;
  wire n30678_o;
  wire n30679_o;
  wire n30680_o;
  wire n30681_o;
  wire n30682_o;
  wire n30683_o;
  wire n30684_o;
  wire n30685_o;
  wire n30686_o;
  wire n30687_o;
  wire n30688_o;
  wire n30689_o;
  wire n30690_o;
  wire n30691_o;
  wire n30692_o;
  wire n30693_o;
  wire n30694_o;
  wire n30695_o;
  wire n30696_o;
  wire n30697_o;
  wire n30698_o;
  wire n30699_o;
  wire n30700_o;
  wire n30701_o;
  wire n30702_o;
  wire n30703_o;
  wire n30704_o;
  wire n30705_o;
  wire n30706_o;
  wire n30707_o;
  wire n30708_o;
  wire n30709_o;
  wire n30710_o;
  wire n30711_o;
  wire n30712_o;
  wire n30713_o;
  wire n30714_o;
  wire n30715_o;
  wire n30716_o;
  wire n30717_o;
  wire n30718_o;
  wire n30719_o;
  wire n30720_o;
  wire n30721_o;
  wire n30722_o;
  wire n30723_o;
  wire n30724_o;
  wire n30725_o;
  wire n30726_o;
  wire [1:0] n30727_o;
  reg n30728_o;
  wire [1:0] n30729_o;
  reg n30730_o;
  wire [1:0] n30731_o;
  reg n30732_o;
  wire [1:0] n30733_o;
  reg n30734_o;
  wire [1:0] n30735_o;
  reg n30736_o;
  wire [1:0] n30737_o;
  reg n30738_o;
  wire [1:0] n30739_o;
  reg n30740_o;
  wire [1:0] n30741_o;
  reg n30742_o;
  wire [1:0] n30743_o;
  reg n30744_o;
  wire [1:0] n30745_o;
  reg n30746_o;
  wire [1:0] n30747_o;
  reg n30748_o;
  wire [1:0] n30749_o;
  reg n30750_o;
  wire [1:0] n30751_o;
  reg n30752_o;
  wire [1:0] n30753_o;
  reg n30754_o;
  wire [1:0] n30755_o;
  reg n30756_o;
  wire [1:0] n30757_o;
  reg n30758_o;
  wire [1:0] n30759_o;
  reg n30760_o;
  wire [1:0] n30761_o;
  reg n30762_o;
  wire [1:0] n30763_o;
  reg n30764_o;
  wire [1:0] n30765_o;
  reg n30766_o;
  wire [1:0] n30767_o;
  reg n30768_o;
  wire n30769_o;
  wire n30770_o;
  wire n30771_o;
  wire n30772_o;
  wire n30773_o;
  wire n30774_o;
  wire n30775_o;
  wire n30776_o;
  wire n30777_o;
  wire n30778_o;
  wire n30779_o;
  wire n30780_o;
  wire n30781_o;
  wire n30782_o;
  wire n30783_o;
  wire n30784_o;
  wire n30785_o;
  wire n30786_o;
  wire n30787_o;
  wire n30788_o;
  wire n30789_o;
  wire n30790_o;
  wire n30791_o;
  wire n30792_o;
  wire n30793_o;
  wire n30794_o;
  wire n30795_o;
  wire n30796_o;
  wire n30797_o;
  wire n30798_o;
  wire n30799_o;
  wire n30800_o;
  wire n30801_o;
  wire n30802_o;
  wire n30803_o;
  wire n30804_o;
  wire n30805_o;
  wire n30806_o;
  wire n30807_o;
  wire n30808_o;
  wire n30809_o;
  wire n30810_o;
  wire n30811_o;
  wire n30812_o;
  wire n30813_o;
  wire n30814_o;
  wire n30815_o;
  wire n30816_o;
  wire n30817_o;
  wire n30818_o;
  wire n30819_o;
  wire n30820_o;
  wire n30821_o;
  wire n30822_o;
  wire n30823_o;
  wire n30824_o;
  wire n30825_o;
  wire n30826_o;
  wire n30827_o;
  wire n30828_o;
  wire n30829_o;
  wire n30830_o;
  wire n30831_o;
  wire n30832_o;
  wire [1:0] n30833_o;
  reg n30834_o;
  wire [1:0] n30835_o;
  reg n30836_o;
  wire [1:0] n30837_o;
  reg n30838_o;
  wire [1:0] n30839_o;
  reg n30840_o;
  wire [1:0] n30841_o;
  reg n30842_o;
  wire [1:0] n30843_o;
  reg n30844_o;
  wire [1:0] n30845_o;
  reg n30846_o;
  wire [1:0] n30847_o;
  reg n30848_o;
  wire [1:0] n30849_o;
  reg n30850_o;
  wire [1:0] n30851_o;
  reg n30852_o;
  wire [1:0] n30853_o;
  reg n30854_o;
  wire [1:0] n30855_o;
  reg n30856_o;
  wire [1:0] n30857_o;
  reg n30858_o;
  wire [1:0] n30859_o;
  reg n30860_o;
  wire [1:0] n30861_o;
  reg n30862_o;
  wire [1:0] n30863_o;
  reg n30864_o;
  wire [1:0] n30865_o;
  reg n30866_o;
  wire [1:0] n30867_o;
  reg n30868_o;
  wire [1:0] n30869_o;
  reg n30870_o;
  wire [1:0] n30871_o;
  reg n30872_o;
  wire [1:0] n30873_o;
  reg n30874_o;
  wire n30875_o;
  wire n30876_o;
  wire n30877_o;
  wire n30878_o;
  wire n30879_o;
  wire n30880_o;
  wire n30881_o;
  wire n30882_o;
  wire n30883_o;
  wire n30884_o;
  wire n30885_o;
  wire n30886_o;
  wire n30887_o;
  wire n30888_o;
  wire n30889_o;
  wire n30890_o;
  wire n30891_o;
  wire n30892_o;
  wire n30893_o;
  wire n30894_o;
  wire n30895_o;
  wire n30896_o;
  wire n30897_o;
  wire n30898_o;
  wire n30899_o;
  wire n30900_o;
  wire n30901_o;
  wire n30902_o;
  wire n30903_o;
  wire n30904_o;
  wire n30905_o;
  wire n30906_o;
  wire n30907_o;
  wire n30908_o;
  wire n30909_o;
  wire n30910_o;
  wire n30911_o;
  wire n30912_o;
  wire n30913_o;
  wire n30914_o;
  wire n30915_o;
  wire n30916_o;
  wire n30917_o;
  wire n30918_o;
  wire n30919_o;
  wire n30920_o;
  wire n30921_o;
  wire n30922_o;
  wire n30923_o;
  wire n30924_o;
  wire n30925_o;
  wire n30926_o;
  wire n30927_o;
  wire n30928_o;
  wire n30929_o;
  wire n30930_o;
  wire n30931_o;
  wire n30932_o;
  wire n30933_o;
  wire n30934_o;
  wire n30935_o;
  wire n30936_o;
  wire n30937_o;
  wire n30938_o;
  wire [1:0] n30939_o;
  reg n30940_o;
  wire [1:0] n30941_o;
  reg n30942_o;
  wire [1:0] n30943_o;
  reg n30944_o;
  wire [1:0] n30945_o;
  reg n30946_o;
  wire [1:0] n30947_o;
  reg n30948_o;
  wire [1:0] n30949_o;
  reg n30950_o;
  wire [1:0] n30951_o;
  reg n30952_o;
  wire [1:0] n30953_o;
  reg n30954_o;
  wire [1:0] n30955_o;
  reg n30956_o;
  wire [1:0] n30957_o;
  reg n30958_o;
  wire [1:0] n30959_o;
  reg n30960_o;
  wire [1:0] n30961_o;
  reg n30962_o;
  wire [1:0] n30963_o;
  reg n30964_o;
  wire [1:0] n30965_o;
  reg n30966_o;
  wire [1:0] n30967_o;
  reg n30968_o;
  wire [1:0] n30969_o;
  reg n30970_o;
  wire [1:0] n30971_o;
  reg n30972_o;
  wire [1:0] n30973_o;
  reg n30974_o;
  wire [1:0] n30975_o;
  reg n30976_o;
  wire [1:0] n30977_o;
  reg n30978_o;
  wire [1:0] n30979_o;
  reg n30980_o;
  wire n30981_o;
  wire n30982_o;
  wire n30983_o;
  wire n30984_o;
  wire n30985_o;
  wire n30986_o;
  wire n30987_o;
  wire n30988_o;
  wire n30989_o;
  wire n30990_o;
  wire n30991_o;
  wire n30992_o;
  wire n30993_o;
  wire n30994_o;
  wire n30995_o;
  wire n30996_o;
  wire n30997_o;
  wire n30998_o;
  wire n30999_o;
  wire n31000_o;
  wire n31001_o;
  wire n31002_o;
  wire n31003_o;
  wire n31004_o;
  wire n31005_o;
  wire n31006_o;
  wire n31007_o;
  wire n31008_o;
  wire n31009_o;
  wire n31010_o;
  wire n31011_o;
  wire n31012_o;
  wire n31013_o;
  wire n31014_o;
  wire n31015_o;
  wire n31016_o;
  wire n31017_o;
  wire n31018_o;
  wire n31019_o;
  wire n31020_o;
  wire n31021_o;
  wire n31022_o;
  wire n31023_o;
  wire n31024_o;
  wire n31025_o;
  wire n31026_o;
  wire n31027_o;
  wire n31028_o;
  wire n31029_o;
  wire n31030_o;
  wire n31031_o;
  wire n31032_o;
  wire n31033_o;
  wire n31034_o;
  wire n31035_o;
  wire n31036_o;
  wire n31037_o;
  wire n31038_o;
  wire n31039_o;
  wire n31040_o;
  wire n31041_o;
  wire n31042_o;
  wire n31043_o;
  wire n31044_o;
  wire [1:0] n31045_o;
  reg n31046_o;
  wire [1:0] n31047_o;
  reg n31048_o;
  wire [1:0] n31049_o;
  reg n31050_o;
  wire [1:0] n31051_o;
  reg n31052_o;
  wire [1:0] n31053_o;
  reg n31054_o;
  wire [1:0] n31055_o;
  reg n31056_o;
  wire [1:0] n31057_o;
  reg n31058_o;
  wire [1:0] n31059_o;
  reg n31060_o;
  wire [1:0] n31061_o;
  reg n31062_o;
  wire [1:0] n31063_o;
  reg n31064_o;
  wire [1:0] n31065_o;
  reg n31066_o;
  wire [1:0] n31067_o;
  reg n31068_o;
  wire [1:0] n31069_o;
  reg n31070_o;
  wire [1:0] n31071_o;
  reg n31072_o;
  wire [1:0] n31073_o;
  reg n31074_o;
  wire [1:0] n31075_o;
  reg n31076_o;
  wire [1:0] n31077_o;
  reg n31078_o;
  wire [1:0] n31079_o;
  reg n31080_o;
  wire [1:0] n31081_o;
  reg n31082_o;
  wire [1:0] n31083_o;
  reg n31084_o;
  wire [1:0] n31085_o;
  reg n31086_o;
  wire n31087_o;
  wire n31088_o;
  wire n31089_o;
  wire n31090_o;
  wire n31091_o;
  wire n31092_o;
  wire n31093_o;
  wire n31094_o;
  wire n31095_o;
  wire n31096_o;
  wire n31097_o;
  wire n31098_o;
  wire n31099_o;
  wire n31100_o;
  wire n31101_o;
  wire n31102_o;
  wire n31103_o;
  wire n31104_o;
  wire n31105_o;
  wire n31106_o;
  wire n31107_o;
  wire n31108_o;
  wire n31109_o;
  wire n31110_o;
  wire n31111_o;
  wire n31112_o;
  wire n31113_o;
  wire n31114_o;
  wire n31115_o;
  wire n31116_o;
  wire n31117_o;
  wire n31118_o;
  wire n31119_o;
  wire n31120_o;
  wire n31121_o;
  wire n31122_o;
  wire n31123_o;
  wire n31124_o;
  wire n31125_o;
  wire n31126_o;
  wire n31127_o;
  wire n31128_o;
  wire n31129_o;
  wire n31130_o;
  wire n31131_o;
  wire n31132_o;
  wire n31133_o;
  wire n31134_o;
  wire n31135_o;
  wire n31136_o;
  wire n31137_o;
  wire n31138_o;
  wire n31139_o;
  wire n31140_o;
  wire n31141_o;
  wire n31142_o;
  wire n31143_o;
  wire n31144_o;
  wire n31145_o;
  wire n31146_o;
  wire n31147_o;
  wire n31148_o;
  wire n31149_o;
  wire n31150_o;
  wire [1:0] n31151_o;
  reg n31152_o;
  wire [1:0] n31153_o;
  reg n31154_o;
  wire [1:0] n31155_o;
  reg n31156_o;
  wire [1:0] n31157_o;
  reg n31158_o;
  wire [1:0] n31159_o;
  reg n31160_o;
  wire [1:0] n31161_o;
  reg n31162_o;
  wire [1:0] n31163_o;
  reg n31164_o;
  wire [1:0] n31165_o;
  reg n31166_o;
  wire [1:0] n31167_o;
  reg n31168_o;
  wire [1:0] n31169_o;
  reg n31170_o;
  wire [1:0] n31171_o;
  reg n31172_o;
  wire [1:0] n31173_o;
  reg n31174_o;
  wire [1:0] n31175_o;
  reg n31176_o;
  wire [1:0] n31177_o;
  reg n31178_o;
  wire [1:0] n31179_o;
  reg n31180_o;
  wire [1:0] n31181_o;
  reg n31182_o;
  wire [1:0] n31183_o;
  reg n31184_o;
  wire [1:0] n31185_o;
  reg n31186_o;
  wire [1:0] n31187_o;
  reg n31188_o;
  wire [1:0] n31189_o;
  reg n31190_o;
  wire [1:0] n31191_o;
  reg n31192_o;
  wire n31193_o;
  wire n31194_o;
  wire n31195_o;
  wire n31196_o;
  wire n31197_o;
  wire n31198_o;
  wire n31199_o;
  wire n31200_o;
  wire n31201_o;
  wire n31202_o;
  wire n31203_o;
  wire n31204_o;
  wire n31205_o;
  wire n31206_o;
  wire n31207_o;
  wire n31208_o;
  wire n31209_o;
  wire n31210_o;
  wire n31211_o;
  wire n31212_o;
  wire n31213_o;
  wire n31214_o;
  wire n31215_o;
  wire n31216_o;
  wire n31217_o;
  wire n31218_o;
  wire n31219_o;
  wire n31220_o;
  wire n31221_o;
  wire n31222_o;
  wire n31223_o;
  wire n31224_o;
  wire n31225_o;
  wire n31226_o;
  wire n31227_o;
  wire n31228_o;
  wire n31229_o;
  wire n31230_o;
  wire n31231_o;
  wire n31232_o;
  wire n31233_o;
  wire n31234_o;
  wire n31235_o;
  wire n31236_o;
  wire n31237_o;
  wire n31238_o;
  wire n31239_o;
  wire n31240_o;
  wire n31241_o;
  wire n31242_o;
  wire n31243_o;
  wire n31244_o;
  wire n31245_o;
  wire n31246_o;
  wire n31247_o;
  wire n31248_o;
  wire n31249_o;
  wire n31250_o;
  wire n31251_o;
  wire n31252_o;
  wire n31253_o;
  wire n31254_o;
  wire n31255_o;
  wire n31256_o;
  wire [1:0] n31257_o;
  reg n31258_o;
  wire [1:0] n31259_o;
  reg n31260_o;
  wire [1:0] n31261_o;
  reg n31262_o;
  wire [1:0] n31263_o;
  reg n31264_o;
  wire [1:0] n31265_o;
  reg n31266_o;
  wire [1:0] n31267_o;
  reg n31268_o;
  wire [1:0] n31269_o;
  reg n31270_o;
  wire [1:0] n31271_o;
  reg n31272_o;
  wire [1:0] n31273_o;
  reg n31274_o;
  wire [1:0] n31275_o;
  reg n31276_o;
  wire [1:0] n31277_o;
  reg n31278_o;
  wire [1:0] n31279_o;
  reg n31280_o;
  wire [1:0] n31281_o;
  reg n31282_o;
  wire [1:0] n31283_o;
  reg n31284_o;
  wire [1:0] n31285_o;
  reg n31286_o;
  wire [1:0] n31287_o;
  reg n31288_o;
  wire [1:0] n31289_o;
  reg n31290_o;
  wire [1:0] n31291_o;
  reg n31292_o;
  wire [1:0] n31293_o;
  reg n31294_o;
  wire [1:0] n31295_o;
  reg n31296_o;
  wire [1:0] n31297_o;
  reg n31298_o;
  assign result = n30445_o;
  /* logical.vhdl:23:12  */
  assign par0 = n28923_o; // (signal)
  /* logical.vhdl:23:18  */
  assign par1 = n28930_o; // (signal)
  /* logical.vhdl:24:12  */
  assign parity = n30449_o; // (signal)
  /* logical.vhdl:25:12  */
  assign permute = n30450_o; // (signal)
  /* logical.vhdl:100:19  */
  assign n28917_o = rs[0];
  /* logical.vhdl:100:29  */
  assign n28918_o = rs[8];
  /* logical.vhdl:100:23  */
  assign n28919_o = n28917_o ^ n28918_o;
  /* logical.vhdl:100:39  */
  assign n28920_o = rs[16];
  /* logical.vhdl:100:33  */
  assign n28921_o = n28919_o ^ n28920_o;
  /* logical.vhdl:100:50  */
  assign n28922_o = rs[24];
  /* logical.vhdl:100:44  */
  assign n28923_o = n28921_o ^ n28922_o;
  /* logical.vhdl:101:19  */
  assign n28924_o = rs[32];
  /* logical.vhdl:101:30  */
  assign n28925_o = rs[40];
  /* logical.vhdl:101:24  */
  assign n28926_o = n28924_o ^ n28925_o;
  /* logical.vhdl:101:41  */
  assign n28927_o = rs[48];
  /* logical.vhdl:101:35  */
  assign n28928_o = n28926_o ^ n28927_o;
  /* logical.vhdl:101:52  */
  assign n28929_o = rs[56];
  /* logical.vhdl:101:46  */
  assign n28930_o = n28928_o ^ n28929_o;
  /* logical.vhdl:103:19  */
  assign n28931_o = datalen[3];
  /* logical.vhdl:104:31  */
  assign n28932_o = par0 ^ par1;
  /* logical.vhdl:103:9  */
  assign n28933_o = n28931_o ? n28932_o : par0;
  /* logical.vhdl:103:9  */
  assign n28935_o = n28931_o ? 1'b0 : par1;
  assign n28938_o = n28936_o[63:33];
  assign n28939_o = n28936_o[31:1];
  /* logical.vhdl:113:18  */
  assign n28940_o = rs[7:6];
  /* logical.vhdl:113:35  */
  assign n28942_o = n28940_o == 2'b00;
  /* logical.vhdl:114:60  */
  assign n28943_o = rs[5:0];
  /* logical.vhdl:114:54  */
  assign n28944_o = ~n28943_o;
  /* logical.vhdl:113:13  */
  assign n28949_o = n28942_o ? n30556_o : 1'b0;
  /* logical.vhdl:113:18  */
  assign n28950_o = rs[15:14];
  /* logical.vhdl:113:35  */
  assign n28952_o = n28950_o == 2'b00;
  /* logical.vhdl:114:60  */
  assign n28953_o = rs[13:8];
  /* logical.vhdl:114:54  */
  assign n28954_o = ~n28953_o;
  /* logical.vhdl:113:13  */
  assign n28959_o = n28952_o ? n30662_o : 1'b0;
  /* logical.vhdl:113:18  */
  assign n28960_o = rs[23:22];
  /* logical.vhdl:113:35  */
  assign n28962_o = n28960_o == 2'b00;
  /* logical.vhdl:114:60  */
  assign n28963_o = rs[21:16];
  /* logical.vhdl:114:54  */
  assign n28964_o = ~n28963_o;
  /* logical.vhdl:113:13  */
  assign n28969_o = n28962_o ? n30768_o : 1'b0;
  /* logical.vhdl:113:18  */
  assign n28970_o = rs[31:30];
  /* logical.vhdl:113:35  */
  assign n28972_o = n28970_o == 2'b00;
  /* logical.vhdl:114:60  */
  assign n28973_o = rs[29:24];
  /* logical.vhdl:114:54  */
  assign n28974_o = ~n28973_o;
  /* logical.vhdl:113:13  */
  assign n28979_o = n28972_o ? n30874_o : 1'b0;
  /* logical.vhdl:113:18  */
  assign n28980_o = rs[39:38];
  /* logical.vhdl:113:35  */
  assign n28982_o = n28980_o == 2'b00;
  /* logical.vhdl:114:60  */
  assign n28983_o = rs[37:32];
  /* logical.vhdl:114:54  */
  assign n28984_o = ~n28983_o;
  /* logical.vhdl:113:13  */
  assign n28989_o = n28982_o ? n30980_o : 1'b0;
  /* logical.vhdl:113:18  */
  assign n28990_o = rs[47:46];
  /* logical.vhdl:113:35  */
  assign n28992_o = n28990_o == 2'b00;
  /* logical.vhdl:114:60  */
  assign n28993_o = rs[45:40];
  /* logical.vhdl:114:54  */
  assign n28994_o = ~n28993_o;
  /* logical.vhdl:113:13  */
  assign n28999_o = n28992_o ? n31086_o : 1'b0;
  /* logical.vhdl:113:18  */
  assign n29000_o = rs[55:54];
  /* logical.vhdl:113:35  */
  assign n29002_o = n29000_o == 2'b00;
  /* logical.vhdl:114:60  */
  assign n29003_o = rs[53:48];
  /* logical.vhdl:114:54  */
  assign n29004_o = ~n29003_o;
  /* logical.vhdl:113:13  */
  assign n29009_o = n29002_o ? n31192_o : 1'b0;
  /* logical.vhdl:113:18  */
  assign n29010_o = rs[63:62];
  /* logical.vhdl:113:35  */
  assign n29012_o = n29010_o == 2'b00;
  /* logical.vhdl:114:60  */
  assign n29013_o = rs[61:56];
  /* logical.vhdl:114:54  */
  assign n29014_o = ~n29013_o;
  /* logical.vhdl:113:13  */
  assign n29019_o = n29012_o ? n31298_o : 1'b0;
  /* logical.vhdl:122:23  */
  assign n29020_o = ~rb;
  /* logical.vhdl:121:9  */
  assign n29021_o = invert_in ? n29020_o : rb;
  /* logical.vhdl:129:35  */
  assign n29022_o = rs & n29021_o;
  /* logical.vhdl:128:21  */
  assign n29024_o = op == 6'b000011;
  /* logical.vhdl:131:35  */
  assign n29025_o = rs | n29021_o;
  /* logical.vhdl:130:21  */
  assign n29027_o = op == 6'b101100;
  /* logical.vhdl:133:35  */
  assign n29028_o = rs ^ n29021_o;
  assign n29029_o = {n29027_o, n29024_o};
  /* logical.vhdl:127:17  */
  always @*
    case (n29029_o)
      2'b10: n29030_o = n29025_o;
      2'b01: n29030_o = n29022_o;
      default: n29030_o = n29028_o;
    endcase
  /* logical.vhdl:136:28  */
  assign n29031_o = ~n29030_o;
  /* logical.vhdl:135:17  */
  assign n29032_o = invert_out ? n29031_o : n29030_o;
  /* logical.vhdl:126:13  */
  assign n29034_o = op == 6'b000011;
  /* logical.vhdl:126:25  */
  assign n29036_o = op == 6'b101100;
  /* logical.vhdl:126:25  */
  assign n29037_o = n29034_o | n29036_o;
  /* logical.vhdl:126:33  */
  assign n29039_o = op == 6'b111010;
  /* logical.vhdl:126:33  */
  assign n29040_o = n29037_o | n29039_o;
  /* logical.vhdl:139:13  */
  assign n29042_o = op == 6'b101110;
  /* ppc_fx_insns.vhdl:745:61  */
  assign n29052_o = rs[7:0];
  /* ppc_fx_insns.vhdl:745:79  */
  assign n29053_o = rb[7:0];
  /* helpers.vhdl:126:14  */
  assign n29059_o = n29052_o == n29053_o;
  /* helpers.vhdl:126:9  */
  assign n29062_o = n29059_o ? 8'b11111111 : 8'b00000000;
  /* ppc_fx_insns.vhdl:745:61  */
  assign n29067_o = rs[15:8];
  /* ppc_fx_insns.vhdl:745:79  */
  assign n29068_o = rb[15:8];
  /* helpers.vhdl:126:14  */
  assign n29074_o = n29067_o == n29068_o;
  /* helpers.vhdl:126:9  */
  assign n29077_o = n29074_o ? 8'b11111111 : 8'b00000000;
  /* ppc_fx_insns.vhdl:745:61  */
  assign n29081_o = rs[23:16];
  /* ppc_fx_insns.vhdl:745:79  */
  assign n29082_o = rb[23:16];
  /* helpers.vhdl:126:14  */
  assign n29088_o = n29081_o == n29082_o;
  /* helpers.vhdl:126:9  */
  assign n29091_o = n29088_o ? 8'b11111111 : 8'b00000000;
  /* ppc_fx_insns.vhdl:745:61  */
  assign n29095_o = rs[31:24];
  /* ppc_fx_insns.vhdl:745:79  */
  assign n29096_o = rb[31:24];
  /* helpers.vhdl:126:14  */
  assign n29102_o = n29095_o == n29096_o;
  /* helpers.vhdl:126:9  */
  assign n29105_o = n29102_o ? 8'b11111111 : 8'b00000000;
  /* ppc_fx_insns.vhdl:745:61  */
  assign n29109_o = rs[39:32];
  /* ppc_fx_insns.vhdl:745:79  */
  assign n29110_o = rb[39:32];
  /* helpers.vhdl:126:14  */
  assign n29116_o = n29109_o == n29110_o;
  /* helpers.vhdl:126:9  */
  assign n29119_o = n29116_o ? 8'b11111111 : 8'b00000000;
  /* ppc_fx_insns.vhdl:745:61  */
  assign n29123_o = rs[47:40];
  /* ppc_fx_insns.vhdl:745:79  */
  assign n29124_o = rb[47:40];
  /* helpers.vhdl:126:14  */
  assign n29130_o = n29123_o == n29124_o;
  /* helpers.vhdl:126:9  */
  assign n29133_o = n29130_o ? 8'b11111111 : 8'b00000000;
  /* ppc_fx_insns.vhdl:745:61  */
  assign n29137_o = rs[55:48];
  /* ppc_fx_insns.vhdl:745:79  */
  assign n29138_o = rb[55:48];
  /* helpers.vhdl:126:14  */
  assign n29144_o = n29137_o == n29138_o;
  /* helpers.vhdl:126:9  */
  assign n29147_o = n29144_o ? 8'b11111111 : 8'b00000000;
  /* ppc_fx_insns.vhdl:745:61  */
  assign n29151_o = rs[63:56];
  /* ppc_fx_insns.vhdl:745:79  */
  assign n29152_o = rb[63:56];
  /* helpers.vhdl:126:14  */
  assign n29158_o = n29151_o == n29152_o;
  /* helpers.vhdl:126:9  */
  assign n29161_o = n29158_o ? 8'b11111111 : 8'b00000000;
  assign n29163_o = {n29161_o, n29147_o, n29133_o, n29119_o, n29105_o, n29091_o, n29077_o, n29062_o};
  /* logical.vhdl:141:13  */
  assign n29165_o = op == 6'b001010;
  /* logical.vhdl:144:42  */
  assign n29166_o = {56'b0, permute};  //  uext
  /* logical.vhdl:143:13  */
  assign n29168_o = op == 6'b001000;
  /* logical.vhdl:147:30  */
  assign n29169_o = ~invert_in;
  /* logical.vhdl:149:50  */
  assign n29171_o = rs[55:44];
  /* logical.vhdl:32:17  */
  assign n29189_o = n29171_o[11];
  /* logical.vhdl:33:17  */
  assign n29191_o = n29171_o[10];
  /* logical.vhdl:34:17  */
  assign n29193_o = n29171_o[9];
  /* logical.vhdl:35:17  */
  assign n29195_o = n29171_o[8];
  /* logical.vhdl:36:17  */
  assign n29197_o = n29171_o[7];
  /* logical.vhdl:37:17  */
  assign n29199_o = n29171_o[6];
  /* logical.vhdl:38:17  */
  assign n29201_o = n29171_o[5];
  /* logical.vhdl:39:17  */
  assign n29203_o = n29171_o[4];
  /* logical.vhdl:40:17  */
  assign n29205_o = n29171_o[3];
  /* logical.vhdl:41:17  */
  assign n29207_o = n29171_o[2];
  /* logical.vhdl:42:17  */
  assign n29209_o = n29171_o[1];
  /* logical.vhdl:43:17  */
  assign n29211_o = n29171_o[0];
  /* logical.vhdl:44:22  */
  assign n29213_o = n29199_o & n29189_o;
  /* logical.vhdl:44:28  */
  assign n29214_o = n29213_o & n29205_o;
  /* logical.vhdl:44:38  */
  assign n29215_o = ~n29197_o;
  /* logical.vhdl:44:34  */
  assign n29216_o = n29214_o & n29215_o;
  /* logical.vhdl:44:51  */
  assign n29217_o = n29207_o & n29189_o;
  /* logical.vhdl:44:61  */
  assign n29218_o = ~n29205_o;
  /* logical.vhdl:44:57  */
  assign n29219_o = n29217_o & n29218_o;
  /* logical.vhdl:44:45  */
  assign n29220_o = n29216_o | n29219_o;
  /* logical.vhdl:44:78  */
  assign n29221_o = ~n29189_o;
  /* logical.vhdl:44:74  */
  assign n29222_o = n29191_o & n29221_o;
  /* logical.vhdl:44:68  */
  assign n29223_o = n29220_o | n29222_o;
  /* logical.vhdl:45:22  */
  assign n29226_o = n29201_o & n29189_o;
  /* logical.vhdl:45:28  */
  assign n29227_o = n29226_o & n29205_o;
  /* logical.vhdl:45:38  */
  assign n29228_o = ~n29197_o;
  /* logical.vhdl:45:34  */
  assign n29229_o = n29227_o & n29228_o;
  /* logical.vhdl:45:51  */
  assign n29230_o = n29209_o & n29189_o;
  /* logical.vhdl:45:61  */
  assign n29231_o = ~n29205_o;
  /* logical.vhdl:45:57  */
  assign n29232_o = n29230_o & n29231_o;
  /* logical.vhdl:45:45  */
  assign n29233_o = n29229_o | n29232_o;
  /* logical.vhdl:45:78  */
  assign n29234_o = ~n29189_o;
  /* logical.vhdl:45:74  */
  assign n29235_o = n29193_o & n29234_o;
  /* logical.vhdl:45:68  */
  assign n29236_o = n29233_o | n29235_o;
  /* logical.vhdl:47:26  */
  assign n29239_o = ~n29189_o;
  /* logical.vhdl:47:22  */
  assign n29240_o = n29207_o & n29239_o;
  /* logical.vhdl:47:32  */
  assign n29241_o = n29240_o & n29197_o;
  /* logical.vhdl:47:42  */
  assign n29242_o = ~n29205_o;
  /* logical.vhdl:47:38  */
  assign n29243_o = n29241_o & n29242_o;
  /* logical.vhdl:47:59  */
  assign n29244_o = ~n29205_o;
  /* logical.vhdl:47:55  */
  assign n29245_o = n29199_o & n29244_o;
  /* logical.vhdl:47:69  */
  assign n29246_o = ~n29197_o;
  /* logical.vhdl:47:65  */
  assign n29247_o = n29245_o & n29246_o;
  /* logical.vhdl:47:49  */
  assign n29248_o = n29243_o | n29247_o;
  /* logical.vhdl:48:26  */
  assign n29249_o = ~n29189_o;
  /* logical.vhdl:48:22  */
  assign n29250_o = n29199_o & n29249_o;
  /* logical.vhdl:48:36  */
  assign n29251_o = ~n29197_o;
  /* logical.vhdl:48:32  */
  assign n29252_o = n29250_o & n29251_o;
  /* logical.vhdl:47:76  */
  assign n29253_o = n29248_o | n29252_o;
  /* logical.vhdl:48:49  */
  assign n29254_o = n29197_o & n29205_o;
  /* logical.vhdl:48:43  */
  assign n29255_o = n29253_o | n29254_o;
  /* logical.vhdl:49:26  */
  assign n29257_o = ~n29189_o;
  /* logical.vhdl:49:22  */
  assign n29258_o = n29209_o & n29257_o;
  /* logical.vhdl:49:32  */
  assign n29259_o = n29258_o & n29197_o;
  /* logical.vhdl:49:42  */
  assign n29260_o = ~n29205_o;
  /* logical.vhdl:49:38  */
  assign n29261_o = n29259_o & n29260_o;
  /* logical.vhdl:49:59  */
  assign n29262_o = ~n29205_o;
  /* logical.vhdl:49:55  */
  assign n29263_o = n29201_o & n29262_o;
  /* logical.vhdl:49:69  */
  assign n29264_o = ~n29197_o;
  /* logical.vhdl:49:65  */
  assign n29265_o = n29263_o & n29264_o;
  /* logical.vhdl:49:49  */
  assign n29266_o = n29261_o | n29265_o;
  /* logical.vhdl:50:26  */
  assign n29267_o = ~n29189_o;
  /* logical.vhdl:50:22  */
  assign n29268_o = n29201_o & n29267_o;
  /* logical.vhdl:50:36  */
  assign n29269_o = ~n29197_o;
  /* logical.vhdl:50:32  */
  assign n29270_o = n29268_o & n29269_o;
  /* logical.vhdl:49:76  */
  assign n29271_o = n29266_o | n29270_o;
  /* logical.vhdl:50:49  */
  assign n29272_o = n29189_o & n29205_o;
  /* logical.vhdl:50:43  */
  assign n29273_o = n29271_o | n29272_o;
  /* logical.vhdl:52:21  */
  assign n29276_o = n29189_o | n29197_o;
  /* logical.vhdl:52:26  */
  assign n29277_o = n29276_o | n29205_o;
  /* logical.vhdl:53:20  */
  assign n29279_o = ~n29197_o;
  /* logical.vhdl:53:26  */
  assign n29280_o = n29279_o & n29207_o;
  /* logical.vhdl:53:36  */
  assign n29281_o = ~n29205_o;
  /* logical.vhdl:53:32  */
  assign n29282_o = n29280_o & n29281_o;
  /* logical.vhdl:53:49  */
  assign n29283_o = n29197_o & n29205_o;
  /* logical.vhdl:53:43  */
  assign n29284_o = n29282_o | n29283_o;
  /* logical.vhdl:53:56  */
  assign n29285_o = n29284_o | n29189_o;
  /* logical.vhdl:54:20  */
  assign n29287_o = ~n29189_o;
  /* logical.vhdl:54:26  */
  assign n29288_o = n29287_o & n29209_o;
  /* logical.vhdl:54:36  */
  assign n29289_o = ~n29205_o;
  /* logical.vhdl:54:32  */
  assign n29290_o = n29288_o & n29289_o;
  /* logical.vhdl:54:49  */
  assign n29291_o = n29189_o & n29205_o;
  /* logical.vhdl:54:43  */
  assign n29292_o = n29290_o | n29291_o;
  /* logical.vhdl:54:56  */
  assign n29293_o = n29292_o | n29197_o;
  assign n29295_o = {n29223_o, n29236_o, n29195_o, n29255_o, n29273_o, n29203_o, n29277_o, n29285_o, n29293_o, n29211_o};
  /* logical.vhdl:149:35  */
  assign n29297_o = {12'b000000000000, n29295_o};
  /* logical.vhdl:149:81  */
  assign n29299_o = rs[43:32];
  /* logical.vhdl:32:17  */
  assign n29317_o = n29299_o[11];
  /* logical.vhdl:33:17  */
  assign n29319_o = n29299_o[10];
  /* logical.vhdl:34:17  */
  assign n29321_o = n29299_o[9];
  /* logical.vhdl:35:17  */
  assign n29323_o = n29299_o[8];
  /* logical.vhdl:36:17  */
  assign n29325_o = n29299_o[7];
  /* logical.vhdl:37:17  */
  assign n29327_o = n29299_o[6];
  /* logical.vhdl:38:17  */
  assign n29329_o = n29299_o[5];
  /* logical.vhdl:39:17  */
  assign n29331_o = n29299_o[4];
  /* logical.vhdl:40:17  */
  assign n29333_o = n29299_o[3];
  /* logical.vhdl:41:17  */
  assign n29335_o = n29299_o[2];
  /* logical.vhdl:42:17  */
  assign n29337_o = n29299_o[1];
  /* logical.vhdl:43:17  */
  assign n29339_o = n29299_o[0];
  /* logical.vhdl:44:22  */
  assign n29341_o = n29327_o & n29317_o;
  /* logical.vhdl:44:28  */
  assign n29342_o = n29341_o & n29333_o;
  /* logical.vhdl:44:38  */
  assign n29343_o = ~n29325_o;
  /* logical.vhdl:44:34  */
  assign n29344_o = n29342_o & n29343_o;
  /* logical.vhdl:44:51  */
  assign n29345_o = n29335_o & n29317_o;
  /* logical.vhdl:44:61  */
  assign n29346_o = ~n29333_o;
  /* logical.vhdl:44:57  */
  assign n29347_o = n29345_o & n29346_o;
  /* logical.vhdl:44:45  */
  assign n29348_o = n29344_o | n29347_o;
  /* logical.vhdl:44:78  */
  assign n29349_o = ~n29317_o;
  /* logical.vhdl:44:74  */
  assign n29350_o = n29319_o & n29349_o;
  /* logical.vhdl:44:68  */
  assign n29351_o = n29348_o | n29350_o;
  /* logical.vhdl:45:22  */
  assign n29354_o = n29329_o & n29317_o;
  /* logical.vhdl:45:28  */
  assign n29355_o = n29354_o & n29333_o;
  /* logical.vhdl:45:38  */
  assign n29356_o = ~n29325_o;
  /* logical.vhdl:45:34  */
  assign n29357_o = n29355_o & n29356_o;
  /* logical.vhdl:45:51  */
  assign n29358_o = n29337_o & n29317_o;
  /* logical.vhdl:45:61  */
  assign n29359_o = ~n29333_o;
  /* logical.vhdl:45:57  */
  assign n29360_o = n29358_o & n29359_o;
  /* logical.vhdl:45:45  */
  assign n29361_o = n29357_o | n29360_o;
  /* logical.vhdl:45:78  */
  assign n29362_o = ~n29317_o;
  /* logical.vhdl:45:74  */
  assign n29363_o = n29321_o & n29362_o;
  /* logical.vhdl:45:68  */
  assign n29364_o = n29361_o | n29363_o;
  /* logical.vhdl:47:26  */
  assign n29367_o = ~n29317_o;
  /* logical.vhdl:47:22  */
  assign n29368_o = n29335_o & n29367_o;
  /* logical.vhdl:47:32  */
  assign n29369_o = n29368_o & n29325_o;
  /* logical.vhdl:47:42  */
  assign n29370_o = ~n29333_o;
  /* logical.vhdl:47:38  */
  assign n29371_o = n29369_o & n29370_o;
  /* logical.vhdl:47:59  */
  assign n29372_o = ~n29333_o;
  /* logical.vhdl:47:55  */
  assign n29373_o = n29327_o & n29372_o;
  /* logical.vhdl:47:69  */
  assign n29374_o = ~n29325_o;
  /* logical.vhdl:47:65  */
  assign n29375_o = n29373_o & n29374_o;
  /* logical.vhdl:47:49  */
  assign n29376_o = n29371_o | n29375_o;
  /* logical.vhdl:48:26  */
  assign n29377_o = ~n29317_o;
  /* logical.vhdl:48:22  */
  assign n29378_o = n29327_o & n29377_o;
  /* logical.vhdl:48:36  */
  assign n29379_o = ~n29325_o;
  /* logical.vhdl:48:32  */
  assign n29380_o = n29378_o & n29379_o;
  /* logical.vhdl:47:76  */
  assign n29381_o = n29376_o | n29380_o;
  /* logical.vhdl:48:49  */
  assign n29382_o = n29325_o & n29333_o;
  /* logical.vhdl:48:43  */
  assign n29383_o = n29381_o | n29382_o;
  /* logical.vhdl:49:26  */
  assign n29385_o = ~n29317_o;
  /* logical.vhdl:49:22  */
  assign n29386_o = n29337_o & n29385_o;
  /* logical.vhdl:49:32  */
  assign n29387_o = n29386_o & n29325_o;
  /* logical.vhdl:49:42  */
  assign n29388_o = ~n29333_o;
  /* logical.vhdl:49:38  */
  assign n29389_o = n29387_o & n29388_o;
  /* logical.vhdl:49:59  */
  assign n29390_o = ~n29333_o;
  /* logical.vhdl:49:55  */
  assign n29391_o = n29329_o & n29390_o;
  /* logical.vhdl:49:69  */
  assign n29392_o = ~n29325_o;
  /* logical.vhdl:49:65  */
  assign n29393_o = n29391_o & n29392_o;
  /* logical.vhdl:49:49  */
  assign n29394_o = n29389_o | n29393_o;
  /* logical.vhdl:50:26  */
  assign n29395_o = ~n29317_o;
  /* logical.vhdl:50:22  */
  assign n29396_o = n29329_o & n29395_o;
  /* logical.vhdl:50:36  */
  assign n29397_o = ~n29325_o;
  /* logical.vhdl:50:32  */
  assign n29398_o = n29396_o & n29397_o;
  /* logical.vhdl:49:76  */
  assign n29399_o = n29394_o | n29398_o;
  /* logical.vhdl:50:49  */
  assign n29400_o = n29317_o & n29333_o;
  /* logical.vhdl:50:43  */
  assign n29401_o = n29399_o | n29400_o;
  /* logical.vhdl:52:21  */
  assign n29404_o = n29317_o | n29325_o;
  /* logical.vhdl:52:26  */
  assign n29405_o = n29404_o | n29333_o;
  /* logical.vhdl:53:20  */
  assign n29407_o = ~n29325_o;
  /* logical.vhdl:53:26  */
  assign n29408_o = n29407_o & n29335_o;
  /* logical.vhdl:53:36  */
  assign n29409_o = ~n29333_o;
  /* logical.vhdl:53:32  */
  assign n29410_o = n29408_o & n29409_o;
  /* logical.vhdl:53:49  */
  assign n29411_o = n29325_o & n29333_o;
  /* logical.vhdl:53:43  */
  assign n29412_o = n29410_o | n29411_o;
  /* logical.vhdl:53:56  */
  assign n29413_o = n29412_o | n29317_o;
  /* logical.vhdl:54:20  */
  assign n29415_o = ~n29317_o;
  /* logical.vhdl:54:26  */
  assign n29416_o = n29415_o & n29337_o;
  /* logical.vhdl:54:36  */
  assign n29417_o = ~n29333_o;
  /* logical.vhdl:54:32  */
  assign n29418_o = n29416_o & n29417_o;
  /* logical.vhdl:54:49  */
  assign n29419_o = n29317_o & n29333_o;
  /* logical.vhdl:54:43  */
  assign n29420_o = n29418_o | n29419_o;
  /* logical.vhdl:54:56  */
  assign n29421_o = n29420_o | n29325_o;
  assign n29423_o = {n29351_o, n29364_o, n29323_o, n29383_o, n29401_o, n29331_o, n29405_o, n29413_o, n29421_o, n29339_o};
  /* logical.vhdl:149:66  */
  assign n29424_o = {n29297_o, n29423_o};
  /* logical.vhdl:149:97  */
  assign n29426_o = {n29424_o, 12'b000000000000};
  /* logical.vhdl:150:50  */
  assign n29428_o = rs[23:12];
  /* logical.vhdl:32:17  */
  assign n29446_o = n29428_o[11];
  /* logical.vhdl:33:17  */
  assign n29448_o = n29428_o[10];
  /* logical.vhdl:34:17  */
  assign n29450_o = n29428_o[9];
  /* logical.vhdl:35:17  */
  assign n29452_o = n29428_o[8];
  /* logical.vhdl:36:17  */
  assign n29454_o = n29428_o[7];
  /* logical.vhdl:37:17  */
  assign n29456_o = n29428_o[6];
  /* logical.vhdl:38:17  */
  assign n29458_o = n29428_o[5];
  /* logical.vhdl:39:17  */
  assign n29460_o = n29428_o[4];
  /* logical.vhdl:40:17  */
  assign n29462_o = n29428_o[3];
  /* logical.vhdl:41:17  */
  assign n29464_o = n29428_o[2];
  /* logical.vhdl:42:17  */
  assign n29466_o = n29428_o[1];
  /* logical.vhdl:43:17  */
  assign n29468_o = n29428_o[0];
  /* logical.vhdl:44:22  */
  assign n29470_o = n29456_o & n29446_o;
  /* logical.vhdl:44:28  */
  assign n29471_o = n29470_o & n29462_o;
  /* logical.vhdl:44:38  */
  assign n29472_o = ~n29454_o;
  /* logical.vhdl:44:34  */
  assign n29473_o = n29471_o & n29472_o;
  /* logical.vhdl:44:51  */
  assign n29474_o = n29464_o & n29446_o;
  /* logical.vhdl:44:61  */
  assign n29475_o = ~n29462_o;
  /* logical.vhdl:44:57  */
  assign n29476_o = n29474_o & n29475_o;
  /* logical.vhdl:44:45  */
  assign n29477_o = n29473_o | n29476_o;
  /* logical.vhdl:44:78  */
  assign n29478_o = ~n29446_o;
  /* logical.vhdl:44:74  */
  assign n29479_o = n29448_o & n29478_o;
  /* logical.vhdl:44:68  */
  assign n29480_o = n29477_o | n29479_o;
  /* logical.vhdl:45:22  */
  assign n29483_o = n29458_o & n29446_o;
  /* logical.vhdl:45:28  */
  assign n29484_o = n29483_o & n29462_o;
  /* logical.vhdl:45:38  */
  assign n29485_o = ~n29454_o;
  /* logical.vhdl:45:34  */
  assign n29486_o = n29484_o & n29485_o;
  /* logical.vhdl:45:51  */
  assign n29487_o = n29466_o & n29446_o;
  /* logical.vhdl:45:61  */
  assign n29488_o = ~n29462_o;
  /* logical.vhdl:45:57  */
  assign n29489_o = n29487_o & n29488_o;
  /* logical.vhdl:45:45  */
  assign n29490_o = n29486_o | n29489_o;
  /* logical.vhdl:45:78  */
  assign n29491_o = ~n29446_o;
  /* logical.vhdl:45:74  */
  assign n29492_o = n29450_o & n29491_o;
  /* logical.vhdl:45:68  */
  assign n29493_o = n29490_o | n29492_o;
  /* logical.vhdl:47:26  */
  assign n29496_o = ~n29446_o;
  /* logical.vhdl:47:22  */
  assign n29497_o = n29464_o & n29496_o;
  /* logical.vhdl:47:32  */
  assign n29498_o = n29497_o & n29454_o;
  /* logical.vhdl:47:42  */
  assign n29499_o = ~n29462_o;
  /* logical.vhdl:47:38  */
  assign n29500_o = n29498_o & n29499_o;
  /* logical.vhdl:47:59  */
  assign n29501_o = ~n29462_o;
  /* logical.vhdl:47:55  */
  assign n29502_o = n29456_o & n29501_o;
  /* logical.vhdl:47:69  */
  assign n29503_o = ~n29454_o;
  /* logical.vhdl:47:65  */
  assign n29504_o = n29502_o & n29503_o;
  /* logical.vhdl:47:49  */
  assign n29505_o = n29500_o | n29504_o;
  /* logical.vhdl:48:26  */
  assign n29506_o = ~n29446_o;
  /* logical.vhdl:48:22  */
  assign n29507_o = n29456_o & n29506_o;
  /* logical.vhdl:48:36  */
  assign n29508_o = ~n29454_o;
  /* logical.vhdl:48:32  */
  assign n29509_o = n29507_o & n29508_o;
  /* logical.vhdl:47:76  */
  assign n29510_o = n29505_o | n29509_o;
  /* logical.vhdl:48:49  */
  assign n29511_o = n29454_o & n29462_o;
  /* logical.vhdl:48:43  */
  assign n29512_o = n29510_o | n29511_o;
  /* logical.vhdl:49:26  */
  assign n29514_o = ~n29446_o;
  /* logical.vhdl:49:22  */
  assign n29515_o = n29466_o & n29514_o;
  /* logical.vhdl:49:32  */
  assign n29516_o = n29515_o & n29454_o;
  /* logical.vhdl:49:42  */
  assign n29517_o = ~n29462_o;
  /* logical.vhdl:49:38  */
  assign n29518_o = n29516_o & n29517_o;
  /* logical.vhdl:49:59  */
  assign n29519_o = ~n29462_o;
  /* logical.vhdl:49:55  */
  assign n29520_o = n29458_o & n29519_o;
  /* logical.vhdl:49:69  */
  assign n29521_o = ~n29454_o;
  /* logical.vhdl:49:65  */
  assign n29522_o = n29520_o & n29521_o;
  /* logical.vhdl:49:49  */
  assign n29523_o = n29518_o | n29522_o;
  /* logical.vhdl:50:26  */
  assign n29524_o = ~n29446_o;
  /* logical.vhdl:50:22  */
  assign n29525_o = n29458_o & n29524_o;
  /* logical.vhdl:50:36  */
  assign n29526_o = ~n29454_o;
  /* logical.vhdl:50:32  */
  assign n29527_o = n29525_o & n29526_o;
  /* logical.vhdl:49:76  */
  assign n29528_o = n29523_o | n29527_o;
  /* logical.vhdl:50:49  */
  assign n29529_o = n29446_o & n29462_o;
  /* logical.vhdl:50:43  */
  assign n29530_o = n29528_o | n29529_o;
  /* logical.vhdl:52:21  */
  assign n29533_o = n29446_o | n29454_o;
  /* logical.vhdl:52:26  */
  assign n29534_o = n29533_o | n29462_o;
  /* logical.vhdl:53:20  */
  assign n29536_o = ~n29454_o;
  /* logical.vhdl:53:26  */
  assign n29537_o = n29536_o & n29464_o;
  /* logical.vhdl:53:36  */
  assign n29538_o = ~n29462_o;
  /* logical.vhdl:53:32  */
  assign n29539_o = n29537_o & n29538_o;
  /* logical.vhdl:53:49  */
  assign n29540_o = n29454_o & n29462_o;
  /* logical.vhdl:53:43  */
  assign n29541_o = n29539_o | n29540_o;
  /* logical.vhdl:53:56  */
  assign n29542_o = n29541_o | n29446_o;
  /* logical.vhdl:54:20  */
  assign n29544_o = ~n29446_o;
  /* logical.vhdl:54:26  */
  assign n29545_o = n29544_o & n29466_o;
  /* logical.vhdl:54:36  */
  assign n29546_o = ~n29462_o;
  /* logical.vhdl:54:32  */
  assign n29547_o = n29545_o & n29546_o;
  /* logical.vhdl:54:49  */
  assign n29548_o = n29446_o & n29462_o;
  /* logical.vhdl:54:43  */
  assign n29549_o = n29547_o | n29548_o;
  /* logical.vhdl:54:56  */
  assign n29550_o = n29549_o | n29454_o;
  assign n29552_o = {n29480_o, n29493_o, n29452_o, n29512_o, n29530_o, n29460_o, n29534_o, n29542_o, n29550_o, n29468_o};
  /* logical.vhdl:150:35  */
  assign n29553_o = {n29426_o, n29552_o};
  /* logical.vhdl:150:81  */
  assign n29555_o = rs[11:0];
  /* logical.vhdl:32:17  */
  assign n29573_o = n29555_o[11];
  /* logical.vhdl:33:17  */
  assign n29575_o = n29555_o[10];
  /* logical.vhdl:34:17  */
  assign n29577_o = n29555_o[9];
  /* logical.vhdl:35:17  */
  assign n29579_o = n29555_o[8];
  /* logical.vhdl:36:17  */
  assign n29581_o = n29555_o[7];
  /* logical.vhdl:37:17  */
  assign n29583_o = n29555_o[6];
  /* logical.vhdl:38:17  */
  assign n29585_o = n29555_o[5];
  /* logical.vhdl:39:17  */
  assign n29587_o = n29555_o[4];
  /* logical.vhdl:40:17  */
  assign n29589_o = n29555_o[3];
  /* logical.vhdl:41:17  */
  assign n29591_o = n29555_o[2];
  /* logical.vhdl:42:17  */
  assign n29593_o = n29555_o[1];
  /* logical.vhdl:43:17  */
  assign n29595_o = n29555_o[0];
  /* logical.vhdl:44:22  */
  assign n29597_o = n29583_o & n29573_o;
  /* logical.vhdl:44:28  */
  assign n29598_o = n29597_o & n29589_o;
  /* logical.vhdl:44:38  */
  assign n29599_o = ~n29581_o;
  /* logical.vhdl:44:34  */
  assign n29600_o = n29598_o & n29599_o;
  /* logical.vhdl:44:51  */
  assign n29601_o = n29591_o & n29573_o;
  /* logical.vhdl:44:61  */
  assign n29602_o = ~n29589_o;
  /* logical.vhdl:44:57  */
  assign n29603_o = n29601_o & n29602_o;
  /* logical.vhdl:44:45  */
  assign n29604_o = n29600_o | n29603_o;
  /* logical.vhdl:44:78  */
  assign n29605_o = ~n29573_o;
  /* logical.vhdl:44:74  */
  assign n29606_o = n29575_o & n29605_o;
  /* logical.vhdl:44:68  */
  assign n29607_o = n29604_o | n29606_o;
  /* logical.vhdl:45:22  */
  assign n29610_o = n29585_o & n29573_o;
  /* logical.vhdl:45:28  */
  assign n29611_o = n29610_o & n29589_o;
  /* logical.vhdl:45:38  */
  assign n29612_o = ~n29581_o;
  /* logical.vhdl:45:34  */
  assign n29613_o = n29611_o & n29612_o;
  /* logical.vhdl:45:51  */
  assign n29614_o = n29593_o & n29573_o;
  /* logical.vhdl:45:61  */
  assign n29615_o = ~n29589_o;
  /* logical.vhdl:45:57  */
  assign n29616_o = n29614_o & n29615_o;
  /* logical.vhdl:45:45  */
  assign n29617_o = n29613_o | n29616_o;
  /* logical.vhdl:45:78  */
  assign n29618_o = ~n29573_o;
  /* logical.vhdl:45:74  */
  assign n29619_o = n29577_o & n29618_o;
  /* logical.vhdl:45:68  */
  assign n29620_o = n29617_o | n29619_o;
  /* logical.vhdl:47:26  */
  assign n29623_o = ~n29573_o;
  /* logical.vhdl:47:22  */
  assign n29624_o = n29591_o & n29623_o;
  /* logical.vhdl:47:32  */
  assign n29625_o = n29624_o & n29581_o;
  /* logical.vhdl:47:42  */
  assign n29626_o = ~n29589_o;
  /* logical.vhdl:47:38  */
  assign n29627_o = n29625_o & n29626_o;
  /* logical.vhdl:47:59  */
  assign n29628_o = ~n29589_o;
  /* logical.vhdl:47:55  */
  assign n29629_o = n29583_o & n29628_o;
  /* logical.vhdl:47:69  */
  assign n29630_o = ~n29581_o;
  /* logical.vhdl:47:65  */
  assign n29631_o = n29629_o & n29630_o;
  /* logical.vhdl:47:49  */
  assign n29632_o = n29627_o | n29631_o;
  /* logical.vhdl:48:26  */
  assign n29633_o = ~n29573_o;
  /* logical.vhdl:48:22  */
  assign n29634_o = n29583_o & n29633_o;
  /* logical.vhdl:48:36  */
  assign n29635_o = ~n29581_o;
  /* logical.vhdl:48:32  */
  assign n29636_o = n29634_o & n29635_o;
  /* logical.vhdl:47:76  */
  assign n29637_o = n29632_o | n29636_o;
  /* logical.vhdl:48:49  */
  assign n29638_o = n29581_o & n29589_o;
  /* logical.vhdl:48:43  */
  assign n29639_o = n29637_o | n29638_o;
  /* logical.vhdl:49:26  */
  assign n29641_o = ~n29573_o;
  /* logical.vhdl:49:22  */
  assign n29642_o = n29593_o & n29641_o;
  /* logical.vhdl:49:32  */
  assign n29643_o = n29642_o & n29581_o;
  /* logical.vhdl:49:42  */
  assign n29644_o = ~n29589_o;
  /* logical.vhdl:49:38  */
  assign n29645_o = n29643_o & n29644_o;
  /* logical.vhdl:49:59  */
  assign n29646_o = ~n29589_o;
  /* logical.vhdl:49:55  */
  assign n29647_o = n29585_o & n29646_o;
  /* logical.vhdl:49:69  */
  assign n29648_o = ~n29581_o;
  /* logical.vhdl:49:65  */
  assign n29649_o = n29647_o & n29648_o;
  /* logical.vhdl:49:49  */
  assign n29650_o = n29645_o | n29649_o;
  /* logical.vhdl:50:26  */
  assign n29651_o = ~n29573_o;
  /* logical.vhdl:50:22  */
  assign n29652_o = n29585_o & n29651_o;
  /* logical.vhdl:50:36  */
  assign n29653_o = ~n29581_o;
  /* logical.vhdl:50:32  */
  assign n29654_o = n29652_o & n29653_o;
  /* logical.vhdl:49:76  */
  assign n29655_o = n29650_o | n29654_o;
  /* logical.vhdl:50:49  */
  assign n29656_o = n29573_o & n29589_o;
  /* logical.vhdl:50:43  */
  assign n29657_o = n29655_o | n29656_o;
  /* logical.vhdl:52:21  */
  assign n29660_o = n29573_o | n29581_o;
  /* logical.vhdl:52:26  */
  assign n29661_o = n29660_o | n29589_o;
  /* logical.vhdl:53:20  */
  assign n29663_o = ~n29581_o;
  /* logical.vhdl:53:26  */
  assign n29664_o = n29663_o & n29591_o;
  /* logical.vhdl:53:36  */
  assign n29665_o = ~n29589_o;
  /* logical.vhdl:53:32  */
  assign n29666_o = n29664_o & n29665_o;
  /* logical.vhdl:53:49  */
  assign n29667_o = n29581_o & n29589_o;
  /* logical.vhdl:53:43  */
  assign n29668_o = n29666_o | n29667_o;
  /* logical.vhdl:53:56  */
  assign n29669_o = n29668_o | n29573_o;
  /* logical.vhdl:54:20  */
  assign n29671_o = ~n29573_o;
  /* logical.vhdl:54:26  */
  assign n29672_o = n29671_o & n29593_o;
  /* logical.vhdl:54:36  */
  assign n29673_o = ~n29589_o;
  /* logical.vhdl:54:32  */
  assign n29674_o = n29672_o & n29673_o;
  /* logical.vhdl:54:49  */
  assign n29675_o = n29573_o & n29589_o;
  /* logical.vhdl:54:43  */
  assign n29676_o = n29674_o | n29675_o;
  /* logical.vhdl:54:56  */
  assign n29677_o = n29676_o | n29581_o;
  assign n29679_o = {n29607_o, n29620_o, n29579_o, n29639_o, n29657_o, n29587_o, n29661_o, n29669_o, n29677_o, n29595_o};
  /* logical.vhdl:150:66  */
  assign n29680_o = {n29553_o, n29679_o};
  /* logical.vhdl:153:49  */
  assign n29682_o = rs[51:42];
  /* logical.vhdl:64:17  */
  assign n29698_o = n29682_o[9];
  /* logical.vhdl:65:17  */
  assign n29700_o = n29682_o[8];
  /* logical.vhdl:66:17  */
  assign n29702_o = n29682_o[7];
  /* logical.vhdl:67:17  */
  assign n29704_o = n29682_o[6];
  /* logical.vhdl:68:17  */
  assign n29706_o = n29682_o[5];
  /* logical.vhdl:69:17  */
  assign n29708_o = n29682_o[4];
  /* logical.vhdl:70:17  */
  assign n29710_o = n29682_o[3];
  /* logical.vhdl:71:17  */
  assign n29712_o = n29682_o[2];
  /* logical.vhdl:72:17  */
  assign n29714_o = n29682_o[1];
  /* logical.vhdl:73:17  */
  assign n29716_o = n29682_o[0];
  /* logical.vhdl:74:21  */
  assign n29718_o = ~n29704_o;
  /* logical.vhdl:74:27  */
  assign n29719_o = n29718_o & n29710_o;
  /* logical.vhdl:74:33  */
  assign n29720_o = n29719_o & n29712_o;
  /* logical.vhdl:74:46  */
  assign n29721_o = n29706_o & n29710_o;
  /* logical.vhdl:74:52  */
  assign n29722_o = n29721_o & n29712_o;
  /* logical.vhdl:74:58  */
  assign n29723_o = n29722_o & n29704_o;
  /* logical.vhdl:74:40  */
  assign n29724_o = n29720_o | n29723_o;
  /* logical.vhdl:74:71  */
  assign n29725_o = n29710_o & n29712_o;
  /* logical.vhdl:74:81  */
  assign n29726_o = ~n29714_o;
  /* logical.vhdl:74:77  */
  assign n29727_o = n29725_o & n29726_o;
  /* logical.vhdl:74:65  */
  assign n29728_o = n29724_o | n29727_o;
  /* logical.vhdl:75:23  */
  assign n29731_o = n29698_o & n29704_o;
  /* logical.vhdl:75:29  */
  assign n29732_o = n29731_o & n29714_o;
  /* logical.vhdl:75:39  */
  assign n29733_o = ~n29706_o;
  /* logical.vhdl:75:35  */
  assign n29734_o = n29732_o & n29733_o;
  /* logical.vhdl:75:56  */
  assign n29735_o = ~n29712_o;
  /* logical.vhdl:75:52  */
  assign n29736_o = n29698_o & n29735_o;
  /* logical.vhdl:75:46  */
  assign n29737_o = n29734_o | n29736_o;
  /* logical.vhdl:75:73  */
  assign n29738_o = ~n29710_o;
  /* logical.vhdl:75:69  */
  assign n29739_o = n29698_o & n29738_o;
  /* logical.vhdl:75:63  */
  assign n29740_o = n29737_o | n29739_o;
  /* logical.vhdl:76:23  */
  assign n29742_o = n29700_o & n29704_o;
  /* logical.vhdl:76:29  */
  assign n29743_o = n29742_o & n29714_o;
  /* logical.vhdl:76:39  */
  assign n29744_o = ~n29706_o;
  /* logical.vhdl:76:35  */
  assign n29745_o = n29743_o & n29744_o;
  /* logical.vhdl:76:56  */
  assign n29746_o = ~n29712_o;
  /* logical.vhdl:76:52  */
  assign n29747_o = n29700_o & n29746_o;
  /* logical.vhdl:76:46  */
  assign n29748_o = n29745_o | n29747_o;
  /* logical.vhdl:76:73  */
  assign n29749_o = ~n29710_o;
  /* logical.vhdl:76:69  */
  assign n29750_o = n29700_o & n29749_o;
  /* logical.vhdl:76:63  */
  assign n29751_o = n29748_o | n29750_o;
  /* logical.vhdl:78:27  */
  assign n29754_o = ~n29712_o;
  /* logical.vhdl:78:23  */
  assign n29755_o = n29710_o & n29754_o;
  /* logical.vhdl:78:33  */
  assign n29756_o = n29755_o & n29714_o;
  /* logical.vhdl:78:46  */
  assign n29757_o = n29704_o & n29710_o;
  /* logical.vhdl:78:52  */
  assign n29758_o = n29757_o & n29712_o;
  /* logical.vhdl:78:58  */
  assign n29759_o = n29758_o & n29714_o;
  /* logical.vhdl:78:40  */
  assign n29760_o = n29756_o | n29759_o;
  /* logical.vhdl:78:69  */
  assign n29761_o = ~n29706_o;
  /* logical.vhdl:78:75  */
  assign n29762_o = n29761_o & n29710_o;
  /* logical.vhdl:78:81  */
  assign n29763_o = n29762_o & n29712_o;
  /* logical.vhdl:78:87  */
  assign n29764_o = n29763_o & n29714_o;
  /* logical.vhdl:78:65  */
  assign n29765_o = n29760_o | n29764_o;
  /* logical.vhdl:79:23  */
  assign n29767_o = n29698_o & n29706_o;
  /* logical.vhdl:79:29  */
  assign n29768_o = n29767_o & n29710_o;
  /* logical.vhdl:79:35  */
  assign n29769_o = n29768_o & n29712_o;
  /* logical.vhdl:79:41  */
  assign n29770_o = n29769_o & n29714_o;
  /* logical.vhdl:79:51  */
  assign n29771_o = ~n29704_o;
  /* logical.vhdl:79:47  */
  assign n29772_o = n29770_o & n29771_o;
  /* logical.vhdl:79:68  */
  assign n29773_o = ~n29714_o;
  /* logical.vhdl:79:64  */
  assign n29774_o = n29704_o & n29773_o;
  /* logical.vhdl:79:74  */
  assign n29775_o = n29774_o & n29710_o;
  /* logical.vhdl:79:58  */
  assign n29776_o = n29772_o | n29775_o;
  /* logical.vhdl:80:27  */
  assign n29777_o = ~n29710_o;
  /* logical.vhdl:80:23  */
  assign n29778_o = n29704_o & n29777_o;
  /* logical.vhdl:79:81  */
  assign n29779_o = n29776_o | n29778_o;
  /* logical.vhdl:81:23  */
  assign n29781_o = n29700_o & n29706_o;
  /* logical.vhdl:81:29  */
  assign n29782_o = n29781_o & n29712_o;
  /* logical.vhdl:81:35  */
  assign n29783_o = n29782_o & n29710_o;
  /* logical.vhdl:81:41  */
  assign n29784_o = n29783_o & n29714_o;
  /* logical.vhdl:81:51  */
  assign n29785_o = ~n29704_o;
  /* logical.vhdl:81:47  */
  assign n29786_o = n29784_o & n29785_o;
  /* logical.vhdl:81:68  */
  assign n29787_o = ~n29714_o;
  /* logical.vhdl:81:64  */
  assign n29788_o = n29706_o & n29787_o;
  /* logical.vhdl:81:74  */
  assign n29789_o = n29788_o & n29710_o;
  /* logical.vhdl:81:58  */
  assign n29790_o = n29786_o | n29789_o;
  /* logical.vhdl:82:27  */
  assign n29791_o = ~n29710_o;
  /* logical.vhdl:82:23  */
  assign n29792_o = n29706_o & n29791_o;
  /* logical.vhdl:81:81  */
  assign n29793_o = n29790_o | n29792_o;
  /* logical.vhdl:84:23  */
  assign n29796_o = n29706_o & n29710_o;
  /* logical.vhdl:84:29  */
  assign n29797_o = n29796_o & n29712_o;
  /* logical.vhdl:84:35  */
  assign n29798_o = n29797_o & n29714_o;
  /* logical.vhdl:84:48  */
  assign n29799_o = n29704_o & n29710_o;
  /* logical.vhdl:84:54  */
  assign n29800_o = n29799_o & n29712_o;
  /* logical.vhdl:84:60  */
  assign n29801_o = n29800_o & n29714_o;
  /* logical.vhdl:84:42  */
  assign n29802_o = n29798_o | n29801_o;
  /* logical.vhdl:84:77  */
  assign n29803_o = ~n29712_o;
  /* logical.vhdl:84:73  */
  assign n29804_o = n29710_o & n29803_o;
  /* logical.vhdl:84:87  */
  assign n29805_o = ~n29714_o;
  /* logical.vhdl:84:83  */
  assign n29806_o = n29804_o & n29805_o;
  /* logical.vhdl:84:67  */
  assign n29807_o = n29802_o | n29806_o;
  /* logical.vhdl:85:27  */
  assign n29809_o = ~n29704_o;
  /* logical.vhdl:85:23  */
  assign n29810_o = n29698_o & n29809_o;
  /* logical.vhdl:85:37  */
  assign n29811_o = ~n29706_o;
  /* logical.vhdl:85:33  */
  assign n29812_o = n29810_o & n29811_o;
  /* logical.vhdl:85:43  */
  assign n29813_o = n29812_o & n29712_o;
  /* logical.vhdl:85:49  */
  assign n29814_o = n29813_o & n29710_o;
  /* logical.vhdl:85:62  */
  assign n29815_o = n29704_o & n29710_o;
  /* logical.vhdl:85:72  */
  assign n29816_o = ~n29712_o;
  /* logical.vhdl:85:68  */
  assign n29817_o = n29815_o & n29816_o;
  /* logical.vhdl:85:78  */
  assign n29818_o = n29817_o & n29714_o;
  /* logical.vhdl:85:56  */
  assign n29819_o = n29814_o | n29818_o;
  /* logical.vhdl:86:23  */
  assign n29820_o = n29698_o & n29712_o;
  /* logical.vhdl:86:33  */
  assign n29821_o = ~n29714_o;
  /* logical.vhdl:86:29  */
  assign n29822_o = n29820_o & n29821_o;
  /* logical.vhdl:86:39  */
  assign n29823_o = n29822_o & n29710_o;
  /* logical.vhdl:85:85  */
  assign n29824_o = n29819_o | n29823_o;
  /* logical.vhdl:86:56  */
  assign n29825_o = ~n29710_o;
  /* logical.vhdl:86:52  */
  assign n29826_o = n29712_o & n29825_o;
  /* logical.vhdl:86:46  */
  assign n29827_o = n29824_o | n29826_o;
  /* logical.vhdl:87:27  */
  assign n29829_o = ~n29704_o;
  /* logical.vhdl:87:23  */
  assign n29830_o = n29700_o & n29829_o;
  /* logical.vhdl:87:37  */
  assign n29831_o = ~n29706_o;
  /* logical.vhdl:87:33  */
  assign n29832_o = n29830_o & n29831_o;
  /* logical.vhdl:87:43  */
  assign n29833_o = n29832_o & n29710_o;
  /* logical.vhdl:87:49  */
  assign n29834_o = n29833_o & n29712_o;
  /* logical.vhdl:87:62  */
  assign n29835_o = n29706_o & n29710_o;
  /* logical.vhdl:87:72  */
  assign n29836_o = ~n29712_o;
  /* logical.vhdl:87:68  */
  assign n29837_o = n29835_o & n29836_o;
  /* logical.vhdl:87:78  */
  assign n29838_o = n29837_o & n29714_o;
  /* logical.vhdl:87:56  */
  assign n29839_o = n29834_o | n29838_o;
  /* logical.vhdl:88:23  */
  assign n29840_o = n29700_o & n29710_o;
  /* logical.vhdl:88:29  */
  assign n29841_o = n29840_o & n29712_o;
  /* logical.vhdl:88:39  */
  assign n29842_o = ~n29714_o;
  /* logical.vhdl:88:35  */
  assign n29843_o = n29841_o & n29842_o;
  /* logical.vhdl:87:85  */
  assign n29844_o = n29839_o | n29843_o;
  /* logical.vhdl:88:56  */
  assign n29845_o = ~n29710_o;
  /* logical.vhdl:88:52  */
  assign n29846_o = n29714_o & n29845_o;
  /* logical.vhdl:88:46  */
  assign n29847_o = n29844_o | n29846_o;
  assign n29849_o = {n29728_o, n29740_o, n29751_o, n29702_o, n29765_o, n29779_o, n29793_o, n29708_o, n29807_o, n29827_o, n29847_o, n29716_o};
  /* logical.vhdl:153:34  */
  assign n29851_o = {8'b00000000, n29849_o};
  /* logical.vhdl:153:80  */
  assign n29853_o = rs[41:32];
  /* logical.vhdl:64:17  */
  assign n29869_o = n29853_o[9];
  /* logical.vhdl:65:17  */
  assign n29871_o = n29853_o[8];
  /* logical.vhdl:66:17  */
  assign n29873_o = n29853_o[7];
  /* logical.vhdl:67:17  */
  assign n29875_o = n29853_o[6];
  /* logical.vhdl:68:17  */
  assign n29877_o = n29853_o[5];
  /* logical.vhdl:69:17  */
  assign n29879_o = n29853_o[4];
  /* logical.vhdl:70:17  */
  assign n29881_o = n29853_o[3];
  /* logical.vhdl:71:17  */
  assign n29883_o = n29853_o[2];
  /* logical.vhdl:72:17  */
  assign n29885_o = n29853_o[1];
  /* logical.vhdl:73:17  */
  assign n29887_o = n29853_o[0];
  /* logical.vhdl:74:21  */
  assign n29889_o = ~n29875_o;
  /* logical.vhdl:74:27  */
  assign n29890_o = n29889_o & n29881_o;
  /* logical.vhdl:74:33  */
  assign n29891_o = n29890_o & n29883_o;
  /* logical.vhdl:74:46  */
  assign n29892_o = n29877_o & n29881_o;
  /* logical.vhdl:74:52  */
  assign n29893_o = n29892_o & n29883_o;
  /* logical.vhdl:74:58  */
  assign n29894_o = n29893_o & n29875_o;
  /* logical.vhdl:74:40  */
  assign n29895_o = n29891_o | n29894_o;
  /* logical.vhdl:74:71  */
  assign n29896_o = n29881_o & n29883_o;
  /* logical.vhdl:74:81  */
  assign n29897_o = ~n29885_o;
  /* logical.vhdl:74:77  */
  assign n29898_o = n29896_o & n29897_o;
  /* logical.vhdl:74:65  */
  assign n29899_o = n29895_o | n29898_o;
  /* logical.vhdl:75:23  */
  assign n29902_o = n29869_o & n29875_o;
  /* logical.vhdl:75:29  */
  assign n29903_o = n29902_o & n29885_o;
  /* logical.vhdl:75:39  */
  assign n29904_o = ~n29877_o;
  /* logical.vhdl:75:35  */
  assign n29905_o = n29903_o & n29904_o;
  /* logical.vhdl:75:56  */
  assign n29906_o = ~n29883_o;
  /* logical.vhdl:75:52  */
  assign n29907_o = n29869_o & n29906_o;
  /* logical.vhdl:75:46  */
  assign n29908_o = n29905_o | n29907_o;
  /* logical.vhdl:75:73  */
  assign n29909_o = ~n29881_o;
  /* logical.vhdl:75:69  */
  assign n29910_o = n29869_o & n29909_o;
  /* logical.vhdl:75:63  */
  assign n29911_o = n29908_o | n29910_o;
  /* logical.vhdl:76:23  */
  assign n29913_o = n29871_o & n29875_o;
  /* logical.vhdl:76:29  */
  assign n29914_o = n29913_o & n29885_o;
  /* logical.vhdl:76:39  */
  assign n29915_o = ~n29877_o;
  /* logical.vhdl:76:35  */
  assign n29916_o = n29914_o & n29915_o;
  /* logical.vhdl:76:56  */
  assign n29917_o = ~n29883_o;
  /* logical.vhdl:76:52  */
  assign n29918_o = n29871_o & n29917_o;
  /* logical.vhdl:76:46  */
  assign n29919_o = n29916_o | n29918_o;
  /* logical.vhdl:76:73  */
  assign n29920_o = ~n29881_o;
  /* logical.vhdl:76:69  */
  assign n29921_o = n29871_o & n29920_o;
  /* logical.vhdl:76:63  */
  assign n29922_o = n29919_o | n29921_o;
  /* logical.vhdl:78:27  */
  assign n29925_o = ~n29883_o;
  /* logical.vhdl:78:23  */
  assign n29926_o = n29881_o & n29925_o;
  /* logical.vhdl:78:33  */
  assign n29927_o = n29926_o & n29885_o;
  /* logical.vhdl:78:46  */
  assign n29928_o = n29875_o & n29881_o;
  /* logical.vhdl:78:52  */
  assign n29929_o = n29928_o & n29883_o;
  /* logical.vhdl:78:58  */
  assign n29930_o = n29929_o & n29885_o;
  /* logical.vhdl:78:40  */
  assign n29931_o = n29927_o | n29930_o;
  /* logical.vhdl:78:69  */
  assign n29932_o = ~n29877_o;
  /* logical.vhdl:78:75  */
  assign n29933_o = n29932_o & n29881_o;
  /* logical.vhdl:78:81  */
  assign n29934_o = n29933_o & n29883_o;
  /* logical.vhdl:78:87  */
  assign n29935_o = n29934_o & n29885_o;
  /* logical.vhdl:78:65  */
  assign n29936_o = n29931_o | n29935_o;
  /* logical.vhdl:79:23  */
  assign n29938_o = n29869_o & n29877_o;
  /* logical.vhdl:79:29  */
  assign n29939_o = n29938_o & n29881_o;
  /* logical.vhdl:79:35  */
  assign n29940_o = n29939_o & n29883_o;
  /* logical.vhdl:79:41  */
  assign n29941_o = n29940_o & n29885_o;
  /* logical.vhdl:79:51  */
  assign n29942_o = ~n29875_o;
  /* logical.vhdl:79:47  */
  assign n29943_o = n29941_o & n29942_o;
  /* logical.vhdl:79:68  */
  assign n29944_o = ~n29885_o;
  /* logical.vhdl:79:64  */
  assign n29945_o = n29875_o & n29944_o;
  /* logical.vhdl:79:74  */
  assign n29946_o = n29945_o & n29881_o;
  /* logical.vhdl:79:58  */
  assign n29947_o = n29943_o | n29946_o;
  /* logical.vhdl:80:27  */
  assign n29948_o = ~n29881_o;
  /* logical.vhdl:80:23  */
  assign n29949_o = n29875_o & n29948_o;
  /* logical.vhdl:79:81  */
  assign n29950_o = n29947_o | n29949_o;
  /* logical.vhdl:81:23  */
  assign n29952_o = n29871_o & n29877_o;
  /* logical.vhdl:81:29  */
  assign n29953_o = n29952_o & n29883_o;
  /* logical.vhdl:81:35  */
  assign n29954_o = n29953_o & n29881_o;
  /* logical.vhdl:81:41  */
  assign n29955_o = n29954_o & n29885_o;
  /* logical.vhdl:81:51  */
  assign n29956_o = ~n29875_o;
  /* logical.vhdl:81:47  */
  assign n29957_o = n29955_o & n29956_o;
  /* logical.vhdl:81:68  */
  assign n29958_o = ~n29885_o;
  /* logical.vhdl:81:64  */
  assign n29959_o = n29877_o & n29958_o;
  /* logical.vhdl:81:74  */
  assign n29960_o = n29959_o & n29881_o;
  /* logical.vhdl:81:58  */
  assign n29961_o = n29957_o | n29960_o;
  /* logical.vhdl:82:27  */
  assign n29962_o = ~n29881_o;
  /* logical.vhdl:82:23  */
  assign n29963_o = n29877_o & n29962_o;
  /* logical.vhdl:81:81  */
  assign n29964_o = n29961_o | n29963_o;
  /* logical.vhdl:84:23  */
  assign n29967_o = n29877_o & n29881_o;
  /* logical.vhdl:84:29  */
  assign n29968_o = n29967_o & n29883_o;
  /* logical.vhdl:84:35  */
  assign n29969_o = n29968_o & n29885_o;
  /* logical.vhdl:84:48  */
  assign n29970_o = n29875_o & n29881_o;
  /* logical.vhdl:84:54  */
  assign n29971_o = n29970_o & n29883_o;
  /* logical.vhdl:84:60  */
  assign n29972_o = n29971_o & n29885_o;
  /* logical.vhdl:84:42  */
  assign n29973_o = n29969_o | n29972_o;
  /* logical.vhdl:84:77  */
  assign n29974_o = ~n29883_o;
  /* logical.vhdl:84:73  */
  assign n29975_o = n29881_o & n29974_o;
  /* logical.vhdl:84:87  */
  assign n29976_o = ~n29885_o;
  /* logical.vhdl:84:83  */
  assign n29977_o = n29975_o & n29976_o;
  /* logical.vhdl:84:67  */
  assign n29978_o = n29973_o | n29977_o;
  /* logical.vhdl:85:27  */
  assign n29980_o = ~n29875_o;
  /* logical.vhdl:85:23  */
  assign n29981_o = n29869_o & n29980_o;
  /* logical.vhdl:85:37  */
  assign n29982_o = ~n29877_o;
  /* logical.vhdl:85:33  */
  assign n29983_o = n29981_o & n29982_o;
  /* logical.vhdl:85:43  */
  assign n29984_o = n29983_o & n29883_o;
  /* logical.vhdl:85:49  */
  assign n29985_o = n29984_o & n29881_o;
  /* logical.vhdl:85:62  */
  assign n29986_o = n29875_o & n29881_o;
  /* logical.vhdl:85:72  */
  assign n29987_o = ~n29883_o;
  /* logical.vhdl:85:68  */
  assign n29988_o = n29986_o & n29987_o;
  /* logical.vhdl:85:78  */
  assign n29989_o = n29988_o & n29885_o;
  /* logical.vhdl:85:56  */
  assign n29990_o = n29985_o | n29989_o;
  /* logical.vhdl:86:23  */
  assign n29991_o = n29869_o & n29883_o;
  /* logical.vhdl:86:33  */
  assign n29992_o = ~n29885_o;
  /* logical.vhdl:86:29  */
  assign n29993_o = n29991_o & n29992_o;
  /* logical.vhdl:86:39  */
  assign n29994_o = n29993_o & n29881_o;
  /* logical.vhdl:85:85  */
  assign n29995_o = n29990_o | n29994_o;
  /* logical.vhdl:86:56  */
  assign n29996_o = ~n29881_o;
  /* logical.vhdl:86:52  */
  assign n29997_o = n29883_o & n29996_o;
  /* logical.vhdl:86:46  */
  assign n29998_o = n29995_o | n29997_o;
  /* logical.vhdl:87:27  */
  assign n30000_o = ~n29875_o;
  /* logical.vhdl:87:23  */
  assign n30001_o = n29871_o & n30000_o;
  /* logical.vhdl:87:37  */
  assign n30002_o = ~n29877_o;
  /* logical.vhdl:87:33  */
  assign n30003_o = n30001_o & n30002_o;
  /* logical.vhdl:87:43  */
  assign n30004_o = n30003_o & n29881_o;
  /* logical.vhdl:87:49  */
  assign n30005_o = n30004_o & n29883_o;
  /* logical.vhdl:87:62  */
  assign n30006_o = n29877_o & n29881_o;
  /* logical.vhdl:87:72  */
  assign n30007_o = ~n29883_o;
  /* logical.vhdl:87:68  */
  assign n30008_o = n30006_o & n30007_o;
  /* logical.vhdl:87:78  */
  assign n30009_o = n30008_o & n29885_o;
  /* logical.vhdl:87:56  */
  assign n30010_o = n30005_o | n30009_o;
  /* logical.vhdl:88:23  */
  assign n30011_o = n29871_o & n29881_o;
  /* logical.vhdl:88:29  */
  assign n30012_o = n30011_o & n29883_o;
  /* logical.vhdl:88:39  */
  assign n30013_o = ~n29885_o;
  /* logical.vhdl:88:35  */
  assign n30014_o = n30012_o & n30013_o;
  /* logical.vhdl:87:85  */
  assign n30015_o = n30010_o | n30014_o;
  /* logical.vhdl:88:56  */
  assign n30016_o = ~n29881_o;
  /* logical.vhdl:88:52  */
  assign n30017_o = n29885_o & n30016_o;
  /* logical.vhdl:88:46  */
  assign n30018_o = n30015_o | n30017_o;
  assign n30020_o = {n29899_o, n29911_o, n29922_o, n29873_o, n29936_o, n29950_o, n29964_o, n29879_o, n29978_o, n29998_o, n30018_o, n29887_o};
  /* logical.vhdl:153:65  */
  assign n30021_o = {n29851_o, n30020_o};
  /* logical.vhdl:153:96  */
  assign n30023_o = {n30021_o, 8'b00000000};
  /* logical.vhdl:154:49  */
  assign n30025_o = rs[19:10];
  /* logical.vhdl:64:17  */
  assign n30041_o = n30025_o[9];
  /* logical.vhdl:65:17  */
  assign n30043_o = n30025_o[8];
  /* logical.vhdl:66:17  */
  assign n30045_o = n30025_o[7];
  /* logical.vhdl:67:17  */
  assign n30047_o = n30025_o[6];
  /* logical.vhdl:68:17  */
  assign n30049_o = n30025_o[5];
  /* logical.vhdl:69:17  */
  assign n30051_o = n30025_o[4];
  /* logical.vhdl:70:17  */
  assign n30053_o = n30025_o[3];
  /* logical.vhdl:71:17  */
  assign n30055_o = n30025_o[2];
  /* logical.vhdl:72:17  */
  assign n30057_o = n30025_o[1];
  /* logical.vhdl:73:17  */
  assign n30059_o = n30025_o[0];
  /* logical.vhdl:74:21  */
  assign n30061_o = ~n30047_o;
  /* logical.vhdl:74:27  */
  assign n30062_o = n30061_o & n30053_o;
  /* logical.vhdl:74:33  */
  assign n30063_o = n30062_o & n30055_o;
  /* logical.vhdl:74:46  */
  assign n30064_o = n30049_o & n30053_o;
  /* logical.vhdl:74:52  */
  assign n30065_o = n30064_o & n30055_o;
  /* logical.vhdl:74:58  */
  assign n30066_o = n30065_o & n30047_o;
  /* logical.vhdl:74:40  */
  assign n30067_o = n30063_o | n30066_o;
  /* logical.vhdl:74:71  */
  assign n30068_o = n30053_o & n30055_o;
  /* logical.vhdl:74:81  */
  assign n30069_o = ~n30057_o;
  /* logical.vhdl:74:77  */
  assign n30070_o = n30068_o & n30069_o;
  /* logical.vhdl:74:65  */
  assign n30071_o = n30067_o | n30070_o;
  /* logical.vhdl:75:23  */
  assign n30074_o = n30041_o & n30047_o;
  /* logical.vhdl:75:29  */
  assign n30075_o = n30074_o & n30057_o;
  /* logical.vhdl:75:39  */
  assign n30076_o = ~n30049_o;
  /* logical.vhdl:75:35  */
  assign n30077_o = n30075_o & n30076_o;
  /* logical.vhdl:75:56  */
  assign n30078_o = ~n30055_o;
  /* logical.vhdl:75:52  */
  assign n30079_o = n30041_o & n30078_o;
  /* logical.vhdl:75:46  */
  assign n30080_o = n30077_o | n30079_o;
  /* logical.vhdl:75:73  */
  assign n30081_o = ~n30053_o;
  /* logical.vhdl:75:69  */
  assign n30082_o = n30041_o & n30081_o;
  /* logical.vhdl:75:63  */
  assign n30083_o = n30080_o | n30082_o;
  /* logical.vhdl:76:23  */
  assign n30085_o = n30043_o & n30047_o;
  /* logical.vhdl:76:29  */
  assign n30086_o = n30085_o & n30057_o;
  /* logical.vhdl:76:39  */
  assign n30087_o = ~n30049_o;
  /* logical.vhdl:76:35  */
  assign n30088_o = n30086_o & n30087_o;
  /* logical.vhdl:76:56  */
  assign n30089_o = ~n30055_o;
  /* logical.vhdl:76:52  */
  assign n30090_o = n30043_o & n30089_o;
  /* logical.vhdl:76:46  */
  assign n30091_o = n30088_o | n30090_o;
  /* logical.vhdl:76:73  */
  assign n30092_o = ~n30053_o;
  /* logical.vhdl:76:69  */
  assign n30093_o = n30043_o & n30092_o;
  /* logical.vhdl:76:63  */
  assign n30094_o = n30091_o | n30093_o;
  /* logical.vhdl:78:27  */
  assign n30097_o = ~n30055_o;
  /* logical.vhdl:78:23  */
  assign n30098_o = n30053_o & n30097_o;
  /* logical.vhdl:78:33  */
  assign n30099_o = n30098_o & n30057_o;
  /* logical.vhdl:78:46  */
  assign n30100_o = n30047_o & n30053_o;
  /* logical.vhdl:78:52  */
  assign n30101_o = n30100_o & n30055_o;
  /* logical.vhdl:78:58  */
  assign n30102_o = n30101_o & n30057_o;
  /* logical.vhdl:78:40  */
  assign n30103_o = n30099_o | n30102_o;
  /* logical.vhdl:78:69  */
  assign n30104_o = ~n30049_o;
  /* logical.vhdl:78:75  */
  assign n30105_o = n30104_o & n30053_o;
  /* logical.vhdl:78:81  */
  assign n30106_o = n30105_o & n30055_o;
  /* logical.vhdl:78:87  */
  assign n30107_o = n30106_o & n30057_o;
  /* logical.vhdl:78:65  */
  assign n30108_o = n30103_o | n30107_o;
  /* logical.vhdl:79:23  */
  assign n30110_o = n30041_o & n30049_o;
  /* logical.vhdl:79:29  */
  assign n30111_o = n30110_o & n30053_o;
  /* logical.vhdl:79:35  */
  assign n30112_o = n30111_o & n30055_o;
  /* logical.vhdl:79:41  */
  assign n30113_o = n30112_o & n30057_o;
  /* logical.vhdl:79:51  */
  assign n30114_o = ~n30047_o;
  /* logical.vhdl:79:47  */
  assign n30115_o = n30113_o & n30114_o;
  /* logical.vhdl:79:68  */
  assign n30116_o = ~n30057_o;
  /* logical.vhdl:79:64  */
  assign n30117_o = n30047_o & n30116_o;
  /* logical.vhdl:79:74  */
  assign n30118_o = n30117_o & n30053_o;
  /* logical.vhdl:79:58  */
  assign n30119_o = n30115_o | n30118_o;
  /* logical.vhdl:80:27  */
  assign n30120_o = ~n30053_o;
  /* logical.vhdl:80:23  */
  assign n30121_o = n30047_o & n30120_o;
  /* logical.vhdl:79:81  */
  assign n30122_o = n30119_o | n30121_o;
  /* logical.vhdl:81:23  */
  assign n30124_o = n30043_o & n30049_o;
  /* logical.vhdl:81:29  */
  assign n30125_o = n30124_o & n30055_o;
  /* logical.vhdl:81:35  */
  assign n30126_o = n30125_o & n30053_o;
  /* logical.vhdl:81:41  */
  assign n30127_o = n30126_o & n30057_o;
  /* logical.vhdl:81:51  */
  assign n30128_o = ~n30047_o;
  /* logical.vhdl:81:47  */
  assign n30129_o = n30127_o & n30128_o;
  /* logical.vhdl:81:68  */
  assign n30130_o = ~n30057_o;
  /* logical.vhdl:81:64  */
  assign n30131_o = n30049_o & n30130_o;
  /* logical.vhdl:81:74  */
  assign n30132_o = n30131_o & n30053_o;
  /* logical.vhdl:81:58  */
  assign n30133_o = n30129_o | n30132_o;
  /* logical.vhdl:82:27  */
  assign n30134_o = ~n30053_o;
  /* logical.vhdl:82:23  */
  assign n30135_o = n30049_o & n30134_o;
  /* logical.vhdl:81:81  */
  assign n30136_o = n30133_o | n30135_o;
  /* logical.vhdl:84:23  */
  assign n30139_o = n30049_o & n30053_o;
  /* logical.vhdl:84:29  */
  assign n30140_o = n30139_o & n30055_o;
  /* logical.vhdl:84:35  */
  assign n30141_o = n30140_o & n30057_o;
  /* logical.vhdl:84:48  */
  assign n30142_o = n30047_o & n30053_o;
  /* logical.vhdl:84:54  */
  assign n30143_o = n30142_o & n30055_o;
  /* logical.vhdl:84:60  */
  assign n30144_o = n30143_o & n30057_o;
  /* logical.vhdl:84:42  */
  assign n30145_o = n30141_o | n30144_o;
  /* logical.vhdl:84:77  */
  assign n30146_o = ~n30055_o;
  /* logical.vhdl:84:73  */
  assign n30147_o = n30053_o & n30146_o;
  /* logical.vhdl:84:87  */
  assign n30148_o = ~n30057_o;
  /* logical.vhdl:84:83  */
  assign n30149_o = n30147_o & n30148_o;
  /* logical.vhdl:84:67  */
  assign n30150_o = n30145_o | n30149_o;
  /* logical.vhdl:85:27  */
  assign n30152_o = ~n30047_o;
  /* logical.vhdl:85:23  */
  assign n30153_o = n30041_o & n30152_o;
  /* logical.vhdl:85:37  */
  assign n30154_o = ~n30049_o;
  /* logical.vhdl:85:33  */
  assign n30155_o = n30153_o & n30154_o;
  /* logical.vhdl:85:43  */
  assign n30156_o = n30155_o & n30055_o;
  /* logical.vhdl:85:49  */
  assign n30157_o = n30156_o & n30053_o;
  /* logical.vhdl:85:62  */
  assign n30158_o = n30047_o & n30053_o;
  /* logical.vhdl:85:72  */
  assign n30159_o = ~n30055_o;
  /* logical.vhdl:85:68  */
  assign n30160_o = n30158_o & n30159_o;
  /* logical.vhdl:85:78  */
  assign n30161_o = n30160_o & n30057_o;
  /* logical.vhdl:85:56  */
  assign n30162_o = n30157_o | n30161_o;
  /* logical.vhdl:86:23  */
  assign n30163_o = n30041_o & n30055_o;
  /* logical.vhdl:86:33  */
  assign n30164_o = ~n30057_o;
  /* logical.vhdl:86:29  */
  assign n30165_o = n30163_o & n30164_o;
  /* logical.vhdl:86:39  */
  assign n30166_o = n30165_o & n30053_o;
  /* logical.vhdl:85:85  */
  assign n30167_o = n30162_o | n30166_o;
  /* logical.vhdl:86:56  */
  assign n30168_o = ~n30053_o;
  /* logical.vhdl:86:52  */
  assign n30169_o = n30055_o & n30168_o;
  /* logical.vhdl:86:46  */
  assign n30170_o = n30167_o | n30169_o;
  /* logical.vhdl:87:27  */
  assign n30172_o = ~n30047_o;
  /* logical.vhdl:87:23  */
  assign n30173_o = n30043_o & n30172_o;
  /* logical.vhdl:87:37  */
  assign n30174_o = ~n30049_o;
  /* logical.vhdl:87:33  */
  assign n30175_o = n30173_o & n30174_o;
  /* logical.vhdl:87:43  */
  assign n30176_o = n30175_o & n30053_o;
  /* logical.vhdl:87:49  */
  assign n30177_o = n30176_o & n30055_o;
  /* logical.vhdl:87:62  */
  assign n30178_o = n30049_o & n30053_o;
  /* logical.vhdl:87:72  */
  assign n30179_o = ~n30055_o;
  /* logical.vhdl:87:68  */
  assign n30180_o = n30178_o & n30179_o;
  /* logical.vhdl:87:78  */
  assign n30181_o = n30180_o & n30057_o;
  /* logical.vhdl:87:56  */
  assign n30182_o = n30177_o | n30181_o;
  /* logical.vhdl:88:23  */
  assign n30183_o = n30043_o & n30053_o;
  /* logical.vhdl:88:29  */
  assign n30184_o = n30183_o & n30055_o;
  /* logical.vhdl:88:39  */
  assign n30185_o = ~n30057_o;
  /* logical.vhdl:88:35  */
  assign n30186_o = n30184_o & n30185_o;
  /* logical.vhdl:87:85  */
  assign n30187_o = n30182_o | n30186_o;
  /* logical.vhdl:88:56  */
  assign n30188_o = ~n30053_o;
  /* logical.vhdl:88:52  */
  assign n30189_o = n30057_o & n30188_o;
  /* logical.vhdl:88:46  */
  assign n30190_o = n30187_o | n30189_o;
  assign n30192_o = {n30071_o, n30083_o, n30094_o, n30045_o, n30108_o, n30122_o, n30136_o, n30051_o, n30150_o, n30170_o, n30190_o, n30059_o};
  /* logical.vhdl:154:34  */
  assign n30193_o = {n30023_o, n30192_o};
  /* logical.vhdl:154:80  */
  assign n30195_o = rs[9:0];
  /* logical.vhdl:64:17  */
  assign n30211_o = n30195_o[9];
  /* logical.vhdl:65:17  */
  assign n30213_o = n30195_o[8];
  /* logical.vhdl:66:17  */
  assign n30215_o = n30195_o[7];
  /* logical.vhdl:67:17  */
  assign n30217_o = n30195_o[6];
  /* logical.vhdl:68:17  */
  assign n30219_o = n30195_o[5];
  /* logical.vhdl:69:17  */
  assign n30221_o = n30195_o[4];
  /* logical.vhdl:70:17  */
  assign n30223_o = n30195_o[3];
  /* logical.vhdl:71:17  */
  assign n30225_o = n30195_o[2];
  /* logical.vhdl:72:17  */
  assign n30227_o = n30195_o[1];
  /* logical.vhdl:73:17  */
  assign n30229_o = n30195_o[0];
  /* logical.vhdl:74:21  */
  assign n30231_o = ~n30217_o;
  /* logical.vhdl:74:27  */
  assign n30232_o = n30231_o & n30223_o;
  /* logical.vhdl:74:33  */
  assign n30233_o = n30232_o & n30225_o;
  /* logical.vhdl:74:46  */
  assign n30234_o = n30219_o & n30223_o;
  /* logical.vhdl:74:52  */
  assign n30235_o = n30234_o & n30225_o;
  /* logical.vhdl:74:58  */
  assign n30236_o = n30235_o & n30217_o;
  /* logical.vhdl:74:40  */
  assign n30237_o = n30233_o | n30236_o;
  /* logical.vhdl:74:71  */
  assign n30238_o = n30223_o & n30225_o;
  /* logical.vhdl:74:81  */
  assign n30239_o = ~n30227_o;
  /* logical.vhdl:74:77  */
  assign n30240_o = n30238_o & n30239_o;
  /* logical.vhdl:74:65  */
  assign n30241_o = n30237_o | n30240_o;
  /* logical.vhdl:75:23  */
  assign n30244_o = n30211_o & n30217_o;
  /* logical.vhdl:75:29  */
  assign n30245_o = n30244_o & n30227_o;
  /* logical.vhdl:75:39  */
  assign n30246_o = ~n30219_o;
  /* logical.vhdl:75:35  */
  assign n30247_o = n30245_o & n30246_o;
  /* logical.vhdl:75:56  */
  assign n30248_o = ~n30225_o;
  /* logical.vhdl:75:52  */
  assign n30249_o = n30211_o & n30248_o;
  /* logical.vhdl:75:46  */
  assign n30250_o = n30247_o | n30249_o;
  /* logical.vhdl:75:73  */
  assign n30251_o = ~n30223_o;
  /* logical.vhdl:75:69  */
  assign n30252_o = n30211_o & n30251_o;
  /* logical.vhdl:75:63  */
  assign n30253_o = n30250_o | n30252_o;
  /* logical.vhdl:76:23  */
  assign n30255_o = n30213_o & n30217_o;
  /* logical.vhdl:76:29  */
  assign n30256_o = n30255_o & n30227_o;
  /* logical.vhdl:76:39  */
  assign n30257_o = ~n30219_o;
  /* logical.vhdl:76:35  */
  assign n30258_o = n30256_o & n30257_o;
  /* logical.vhdl:76:56  */
  assign n30259_o = ~n30225_o;
  /* logical.vhdl:76:52  */
  assign n30260_o = n30213_o & n30259_o;
  /* logical.vhdl:76:46  */
  assign n30261_o = n30258_o | n30260_o;
  /* logical.vhdl:76:73  */
  assign n30262_o = ~n30223_o;
  /* logical.vhdl:76:69  */
  assign n30263_o = n30213_o & n30262_o;
  /* logical.vhdl:76:63  */
  assign n30264_o = n30261_o | n30263_o;
  /* logical.vhdl:78:27  */
  assign n30267_o = ~n30225_o;
  /* logical.vhdl:78:23  */
  assign n30268_o = n30223_o & n30267_o;
  /* logical.vhdl:78:33  */
  assign n30269_o = n30268_o & n30227_o;
  /* logical.vhdl:78:46  */
  assign n30270_o = n30217_o & n30223_o;
  /* logical.vhdl:78:52  */
  assign n30271_o = n30270_o & n30225_o;
  /* logical.vhdl:78:58  */
  assign n30272_o = n30271_o & n30227_o;
  /* logical.vhdl:78:40  */
  assign n30273_o = n30269_o | n30272_o;
  /* logical.vhdl:78:69  */
  assign n30274_o = ~n30219_o;
  /* logical.vhdl:78:75  */
  assign n30275_o = n30274_o & n30223_o;
  /* logical.vhdl:78:81  */
  assign n30276_o = n30275_o & n30225_o;
  /* logical.vhdl:78:87  */
  assign n30277_o = n30276_o & n30227_o;
  /* logical.vhdl:78:65  */
  assign n30278_o = n30273_o | n30277_o;
  /* logical.vhdl:79:23  */
  assign n30280_o = n30211_o & n30219_o;
  /* logical.vhdl:79:29  */
  assign n30281_o = n30280_o & n30223_o;
  /* logical.vhdl:79:35  */
  assign n30282_o = n30281_o & n30225_o;
  /* logical.vhdl:79:41  */
  assign n30283_o = n30282_o & n30227_o;
  /* logical.vhdl:79:51  */
  assign n30284_o = ~n30217_o;
  /* logical.vhdl:79:47  */
  assign n30285_o = n30283_o & n30284_o;
  /* logical.vhdl:79:68  */
  assign n30286_o = ~n30227_o;
  /* logical.vhdl:79:64  */
  assign n30287_o = n30217_o & n30286_o;
  /* logical.vhdl:79:74  */
  assign n30288_o = n30287_o & n30223_o;
  /* logical.vhdl:79:58  */
  assign n30289_o = n30285_o | n30288_o;
  /* logical.vhdl:80:27  */
  assign n30290_o = ~n30223_o;
  /* logical.vhdl:80:23  */
  assign n30291_o = n30217_o & n30290_o;
  /* logical.vhdl:79:81  */
  assign n30292_o = n30289_o | n30291_o;
  /* logical.vhdl:81:23  */
  assign n30294_o = n30213_o & n30219_o;
  /* logical.vhdl:81:29  */
  assign n30295_o = n30294_o & n30225_o;
  /* logical.vhdl:81:35  */
  assign n30296_o = n30295_o & n30223_o;
  /* logical.vhdl:81:41  */
  assign n30297_o = n30296_o & n30227_o;
  /* logical.vhdl:81:51  */
  assign n30298_o = ~n30217_o;
  /* logical.vhdl:81:47  */
  assign n30299_o = n30297_o & n30298_o;
  /* logical.vhdl:81:68  */
  assign n30300_o = ~n30227_o;
  /* logical.vhdl:81:64  */
  assign n30301_o = n30219_o & n30300_o;
  /* logical.vhdl:81:74  */
  assign n30302_o = n30301_o & n30223_o;
  /* logical.vhdl:81:58  */
  assign n30303_o = n30299_o | n30302_o;
  /* logical.vhdl:82:27  */
  assign n30304_o = ~n30223_o;
  /* logical.vhdl:82:23  */
  assign n30305_o = n30219_o & n30304_o;
  /* logical.vhdl:81:81  */
  assign n30306_o = n30303_o | n30305_o;
  /* logical.vhdl:84:23  */
  assign n30309_o = n30219_o & n30223_o;
  /* logical.vhdl:84:29  */
  assign n30310_o = n30309_o & n30225_o;
  /* logical.vhdl:84:35  */
  assign n30311_o = n30310_o & n30227_o;
  /* logical.vhdl:84:48  */
  assign n30312_o = n30217_o & n30223_o;
  /* logical.vhdl:84:54  */
  assign n30313_o = n30312_o & n30225_o;
  /* logical.vhdl:84:60  */
  assign n30314_o = n30313_o & n30227_o;
  /* logical.vhdl:84:42  */
  assign n30315_o = n30311_o | n30314_o;
  /* logical.vhdl:84:77  */
  assign n30316_o = ~n30225_o;
  /* logical.vhdl:84:73  */
  assign n30317_o = n30223_o & n30316_o;
  /* logical.vhdl:84:87  */
  assign n30318_o = ~n30227_o;
  /* logical.vhdl:84:83  */
  assign n30319_o = n30317_o & n30318_o;
  /* logical.vhdl:84:67  */
  assign n30320_o = n30315_o | n30319_o;
  /* logical.vhdl:85:27  */
  assign n30322_o = ~n30217_o;
  /* logical.vhdl:85:23  */
  assign n30323_o = n30211_o & n30322_o;
  /* logical.vhdl:85:37  */
  assign n30324_o = ~n30219_o;
  /* logical.vhdl:85:33  */
  assign n30325_o = n30323_o & n30324_o;
  /* logical.vhdl:85:43  */
  assign n30326_o = n30325_o & n30225_o;
  /* logical.vhdl:85:49  */
  assign n30327_o = n30326_o & n30223_o;
  /* logical.vhdl:85:62  */
  assign n30328_o = n30217_o & n30223_o;
  /* logical.vhdl:85:72  */
  assign n30329_o = ~n30225_o;
  /* logical.vhdl:85:68  */
  assign n30330_o = n30328_o & n30329_o;
  /* logical.vhdl:85:78  */
  assign n30331_o = n30330_o & n30227_o;
  /* logical.vhdl:85:56  */
  assign n30332_o = n30327_o | n30331_o;
  /* logical.vhdl:86:23  */
  assign n30333_o = n30211_o & n30225_o;
  /* logical.vhdl:86:33  */
  assign n30334_o = ~n30227_o;
  /* logical.vhdl:86:29  */
  assign n30335_o = n30333_o & n30334_o;
  /* logical.vhdl:86:39  */
  assign n30336_o = n30335_o & n30223_o;
  /* logical.vhdl:85:85  */
  assign n30337_o = n30332_o | n30336_o;
  /* logical.vhdl:86:56  */
  assign n30338_o = ~n30223_o;
  /* logical.vhdl:86:52  */
  assign n30339_o = n30225_o & n30338_o;
  /* logical.vhdl:86:46  */
  assign n30340_o = n30337_o | n30339_o;
  /* logical.vhdl:87:27  */
  assign n30342_o = ~n30217_o;
  /* logical.vhdl:87:23  */
  assign n30343_o = n30213_o & n30342_o;
  /* logical.vhdl:87:37  */
  assign n30344_o = ~n30219_o;
  /* logical.vhdl:87:33  */
  assign n30345_o = n30343_o & n30344_o;
  /* logical.vhdl:87:43  */
  assign n30346_o = n30345_o & n30223_o;
  /* logical.vhdl:87:49  */
  assign n30347_o = n30346_o & n30225_o;
  /* logical.vhdl:87:62  */
  assign n30348_o = n30219_o & n30223_o;
  /* logical.vhdl:87:72  */
  assign n30349_o = ~n30225_o;
  /* logical.vhdl:87:68  */
  assign n30350_o = n30348_o & n30349_o;
  /* logical.vhdl:87:78  */
  assign n30351_o = n30350_o & n30227_o;
  /* logical.vhdl:87:56  */
  assign n30352_o = n30347_o | n30351_o;
  /* logical.vhdl:88:23  */
  assign n30353_o = n30213_o & n30223_o;
  /* logical.vhdl:88:29  */
  assign n30354_o = n30353_o & n30225_o;
  /* logical.vhdl:88:39  */
  assign n30355_o = ~n30227_o;
  /* logical.vhdl:88:35  */
  assign n30356_o = n30354_o & n30355_o;
  /* logical.vhdl:87:85  */
  assign n30357_o = n30352_o | n30356_o;
  /* logical.vhdl:88:56  */
  assign n30358_o = ~n30223_o;
  /* logical.vhdl:88:52  */
  assign n30359_o = n30227_o & n30358_o;
  /* logical.vhdl:88:46  */
  assign n30360_o = n30357_o | n30359_o;
  assign n30362_o = {n30241_o, n30253_o, n30264_o, n30215_o, n30278_o, n30292_o, n30306_o, n30221_o, n30320_o, n30340_o, n30360_o, n30229_o};
  /* logical.vhdl:154:65  */
  assign n30363_o = {n30193_o, n30362_o};
  /* logical.vhdl:147:17  */
  assign n30364_o = n29169_o ? n29680_o : n30363_o;
  /* logical.vhdl:145:13  */
  assign n30366_o = op == 6'b111011;
  /* logical.vhdl:158:37  */
  assign n30367_o = datalen[0];
  /* logical.vhdl:158:47  */
  assign n30368_o = rs[7];
  /* logical.vhdl:158:41  */
  assign n30369_o = n30367_o & n30368_o;
  /* logical.vhdl:159:37  */
  assign n30370_o = datalen[1];
  /* logical.vhdl:159:47  */
  assign n30371_o = rs[15];
  /* logical.vhdl:159:41  */
  assign n30372_o = n30370_o & n30371_o;
  /* logical.vhdl:158:52  */
  assign n30373_o = n30369_o | n30372_o;
  /* logical.vhdl:160:37  */
  assign n30374_o = datalen[2];
  /* logical.vhdl:160:47  */
  assign n30375_o = rs[31];
  /* logical.vhdl:160:41  */
  assign n30376_o = n30374_o & n30375_o;
  /* logical.vhdl:159:53  */
  assign n30377_o = n30373_o | n30376_o;
  assign n30378_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30379_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30380_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30381_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30382_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30383_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30384_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30385_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30386_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30387_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30388_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30389_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30390_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30391_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30392_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30393_o = {n30377_o, n30377_o, n30377_o, n30377_o};
  assign n30394_o = {n30378_o, n30379_o, n30380_o, n30381_o};
  assign n30395_o = {n30382_o, n30383_o, n30384_o, n30385_o};
  assign n30396_o = {n30386_o, n30387_o, n30388_o, n30389_o};
  assign n30397_o = {n30390_o, n30391_o, n30392_o, n30393_o};
  assign n30398_o = {n30394_o, n30395_o, n30396_o, n30397_o};
  /* logical.vhdl:162:27  */
  assign n30399_o = datalen[2];
  /* logical.vhdl:163:44  */
  assign n30400_o = rs[31:16];
  assign n30401_o = n30398_o[31:16];
  /* logical.vhdl:162:17  */
  assign n30402_o = n30399_o ? n30400_o : n30401_o;
  assign n30403_o = n30398_o[63:32];
  /* logical.vhdl:165:27  */
  assign n30405_o = datalen[2];
  /* logical.vhdl:165:47  */
  assign n30406_o = datalen[1];
  /* logical.vhdl:165:37  */
  assign n30407_o = n30405_o | n30406_o;
  /* logical.vhdl:166:43  */
  assign n30408_o = rs[15:8];
  assign n30409_o = n30398_o[15:8];
  /* logical.vhdl:165:17  */
  assign n30410_o = n30407_o ? n30408_o : n30409_o;
  /* logical.vhdl:168:38  */
  assign n30412_o = rs[7:0];
  /* logical.vhdl:156:13  */
  assign n30414_o = op == 6'b010111;
  assign n30415_o = {n30414_o, n30366_o, n29168_o, n29165_o, n29042_o, n29040_o};
  assign n30416_o = n29032_o[7:0];
  assign n30417_o = parity[7:0];
  assign n30418_o = n29163_o[7:0];
  assign n30419_o = n29166_o[7:0];
  assign n30420_o = n30364_o[7:0];
  assign n30421_o = rs[7:0];
  /* logical.vhdl:125:9  */
  always @*
    case (n30415_o)
      6'b100000: n30422_o = n30412_o;
      6'b010000: n30422_o = n30420_o;
      6'b001000: n30422_o = n30419_o;
      6'b000100: n30422_o = n30418_o;
      6'b000010: n30422_o = n30417_o;
      6'b000001: n30422_o = n30416_o;
      default: n30422_o = n30421_o;
    endcase
  assign n30423_o = n29032_o[15:8];
  assign n30424_o = parity[15:8];
  assign n30425_o = n29163_o[15:8];
  assign n30426_o = n29166_o[15:8];
  assign n30427_o = n30364_o[15:8];
  assign n30428_o = rs[15:8];
  /* logical.vhdl:125:9  */
  always @*
    case (n30415_o)
      6'b100000: n30429_o = n30410_o;
      6'b010000: n30429_o = n30427_o;
      6'b001000: n30429_o = n30426_o;
      6'b000100: n30429_o = n30425_o;
      6'b000010: n30429_o = n30424_o;
      6'b000001: n30429_o = n30423_o;
      default: n30429_o = n30428_o;
    endcase
  assign n30430_o = n29032_o[31:16];
  assign n30431_o = parity[31:16];
  assign n30432_o = n29163_o[31:16];
  assign n30433_o = n29166_o[31:16];
  assign n30434_o = n30364_o[31:16];
  assign n30435_o = rs[31:16];
  /* logical.vhdl:125:9  */
  always @*
    case (n30415_o)
      6'b100000: n30436_o = n30402_o;
      6'b010000: n30436_o = n30434_o;
      6'b001000: n30436_o = n30433_o;
      6'b000100: n30436_o = n30432_o;
      6'b000010: n30436_o = n30431_o;
      6'b000001: n30436_o = n30430_o;
      default: n30436_o = n30435_o;
    endcase
  assign n30437_o = n29032_o[63:32];
  assign n30438_o = parity[63:32];
  assign n30439_o = n29163_o[63:32];
  assign n30440_o = n29166_o[63:32];
  assign n30441_o = n30364_o[63:32];
  assign n30442_o = rs[63:32];
  /* logical.vhdl:125:9  */
  always @*
    case (n30415_o)
      6'b100000: n30443_o = n30403_o;
      6'b010000: n30443_o = n30441_o;
      6'b001000: n30443_o = n30440_o;
      6'b000100: n30443_o = n30439_o;
      6'b000010: n30443_o = n30438_o;
      6'b000001: n30443_o = n30437_o;
      default: n30443_o = n30442_o;
    endcase
  assign n30445_o = {n30443_o, n30436_o, n30429_o, n30422_o};
  assign n30449_o = {n28938_o, n28935_o, n28939_o, n28933_o};
  assign n30450_o = {n29019_o, n29009_o, n28999_o, n28989_o, n28979_o, n28969_o, n28959_o, n28949_o};
  /* logical.vhdl:16:9  */
  assign n30451_o = rb[0];
  assign n30452_o = rb[1];
  assign n30453_o = rb[2];
  assign n30454_o = rb[3];
  /* logical.vhdl:125:9  */
  assign n30455_o = rb[4];
  assign n30456_o = rb[5];
  assign n30457_o = rb[6];
  assign n30458_o = rb[7];
  assign n30459_o = rb[8];
  assign n30460_o = rb[9];
  assign n30461_o = rb[10];
  assign n30462_o = rb[11];
  assign n30463_o = rb[12];
  assign n30464_o = rb[13];
  assign n30465_o = rb[14];
  assign n30466_o = rb[15];
  assign n30467_o = rb[16];
  assign n30468_o = rb[17];
  assign n30469_o = rb[18];
  assign n30470_o = rb[19];
  assign n30471_o = rb[20];
  assign n30472_o = rb[21];
  assign n30473_o = rb[22];
  assign n30474_o = rb[23];
  assign n30475_o = rb[24];
  assign n30476_o = rb[25];
  assign n30477_o = rb[26];
  assign n30478_o = rb[27];
  assign n30479_o = rb[28];
  /* logical.vhdl:61:45  */
  assign n30480_o = rb[29];
  assign n30481_o = rb[30];
  /* logical.vhdl:61:42  */
  assign n30482_o = rb[31];
  assign n30483_o = rb[32];
  /* logical.vhdl:61:39  */
  assign n30484_o = rb[33];
  assign n30485_o = rb[34];
  /* logical.vhdl:61:36  */
  assign n30486_o = rb[35];
  assign n30487_o = rb[36];
  /* logical.vhdl:61:33  */
  assign n30488_o = rb[37];
  assign n30489_o = rb[38];
  /* logical.vhdl:61:30  */
  assign n30490_o = rb[39];
  assign n30491_o = rb[40];
  /* logical.vhdl:61:27  */
  assign n30492_o = rb[41];
  assign n30493_o = rb[42];
  /* logical.vhdl:61:24  */
  assign n30494_o = rb[43];
  assign n30495_o = rb[44];
  /* logical.vhdl:61:21  */
  assign n30496_o = rb[45];
  assign n30497_o = rb[46];
  /* logical.vhdl:61:18  */
  assign n30498_o = rb[47];
  assign n30499_o = rb[48];
  /* logical.vhdl:60:18  */
  assign n30500_o = rb[49];
  assign n30501_o = rb[50];
  /* logical.vhdl:59:14  */
  assign n30502_o = rb[51];
  /* logical.vhdl:59:14  */
  assign n30503_o = rb[52];
  assign n30504_o = rb[53];
  /* logical.vhdl:59:14  */
  assign n30505_o = rb[54];
  assign n30506_o = rb[55];
  assign n30507_o = rb[56];
  assign n30508_o = rb[57];
  assign n30509_o = rb[58];
  assign n30510_o = rb[59];
  assign n30511_o = rb[60];
  assign n30512_o = rb[61];
  assign n30513_o = rb[62];
  assign n30514_o = rb[63];
  /* logical.vhdl:114:33  */
  assign n30515_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30515_o)
      2'b00: n30516_o = n30451_o;
      2'b01: n30516_o = n30452_o;
      2'b10: n30516_o = n30453_o;
      2'b11: n30516_o = n30454_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30517_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30517_o)
      2'b00: n30518_o = n30455_o;
      2'b01: n30518_o = n30456_o;
      2'b10: n30518_o = n30457_o;
      2'b11: n30518_o = n30458_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30519_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30519_o)
      2'b00: n30520_o = n30459_o;
      2'b01: n30520_o = n30460_o;
      2'b10: n30520_o = n30461_o;
      2'b11: n30520_o = n30462_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30521_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30521_o)
      2'b00: n30522_o = n30463_o;
      2'b01: n30522_o = n30464_o;
      2'b10: n30522_o = n30465_o;
      2'b11: n30522_o = n30466_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30523_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30523_o)
      2'b00: n30524_o = n30467_o;
      2'b01: n30524_o = n30468_o;
      2'b10: n30524_o = n30469_o;
      2'b11: n30524_o = n30470_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30525_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30525_o)
      2'b00: n30526_o = n30471_o;
      2'b01: n30526_o = n30472_o;
      2'b10: n30526_o = n30473_o;
      2'b11: n30526_o = n30474_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30527_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30527_o)
      2'b00: n30528_o = n30475_o;
      2'b01: n30528_o = n30476_o;
      2'b10: n30528_o = n30477_o;
      2'b11: n30528_o = n30478_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30529_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30529_o)
      2'b00: n30530_o = n30479_o;
      2'b01: n30530_o = n30480_o;
      2'b10: n30530_o = n30481_o;
      2'b11: n30530_o = n30482_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30531_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30531_o)
      2'b00: n30532_o = n30483_o;
      2'b01: n30532_o = n30484_o;
      2'b10: n30532_o = n30485_o;
      2'b11: n30532_o = n30486_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30533_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30533_o)
      2'b00: n30534_o = n30487_o;
      2'b01: n30534_o = n30488_o;
      2'b10: n30534_o = n30489_o;
      2'b11: n30534_o = n30490_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30535_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30535_o)
      2'b00: n30536_o = n30491_o;
      2'b01: n30536_o = n30492_o;
      2'b10: n30536_o = n30493_o;
      2'b11: n30536_o = n30494_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30537_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30537_o)
      2'b00: n30538_o = n30495_o;
      2'b01: n30538_o = n30496_o;
      2'b10: n30538_o = n30497_o;
      2'b11: n30538_o = n30498_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30539_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30539_o)
      2'b00: n30540_o = n30499_o;
      2'b01: n30540_o = n30500_o;
      2'b10: n30540_o = n30501_o;
      2'b11: n30540_o = n30502_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30541_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30541_o)
      2'b00: n30542_o = n30503_o;
      2'b01: n30542_o = n30504_o;
      2'b10: n30542_o = n30505_o;
      2'b11: n30542_o = n30506_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30543_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30543_o)
      2'b00: n30544_o = n30507_o;
      2'b01: n30544_o = n30508_o;
      2'b10: n30544_o = n30509_o;
      2'b11: n30544_o = n30510_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30545_o = n28944_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30545_o)
      2'b00: n30546_o = n30511_o;
      2'b01: n30546_o = n30512_o;
      2'b10: n30546_o = n30513_o;
      2'b11: n30546_o = n30514_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30547_o = n28944_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30547_o)
      2'b00: n30548_o = n30516_o;
      2'b01: n30548_o = n30518_o;
      2'b10: n30548_o = n30520_o;
      2'b11: n30548_o = n30522_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30549_o = n28944_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30549_o)
      2'b00: n30550_o = n30524_o;
      2'b01: n30550_o = n30526_o;
      2'b10: n30550_o = n30528_o;
      2'b11: n30550_o = n30530_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30551_o = n28944_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30551_o)
      2'b00: n30552_o = n30532_o;
      2'b01: n30552_o = n30534_o;
      2'b10: n30552_o = n30536_o;
      2'b11: n30552_o = n30538_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30553_o = n28944_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30553_o)
      2'b00: n30554_o = n30540_o;
      2'b01: n30554_o = n30542_o;
      2'b10: n30554_o = n30544_o;
      2'b11: n30554_o = n30546_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30555_o = n28944_o[5:4];
  /* logical.vhdl:114:33  */
  always @*
    case (n30555_o)
      2'b00: n30556_o = n30548_o;
      2'b01: n30556_o = n30550_o;
      2'b10: n30556_o = n30552_o;
      2'b11: n30556_o = n30554_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30557_o = rb[0];
  /* logical.vhdl:114:34  */
  assign n30558_o = rb[1];
  assign n30559_o = rb[2];
  assign n30560_o = rb[3];
  assign n30561_o = rb[4];
  assign n30562_o = rb[5];
  assign n30563_o = rb[6];
  assign n30564_o = rb[7];
  assign n30565_o = rb[8];
  assign n30566_o = rb[9];
  assign n30567_o = rb[10];
  assign n30568_o = rb[11];
  assign n30569_o = rb[12];
  assign n30570_o = rb[13];
  assign n30571_o = rb[14];
  assign n30572_o = rb[15];
  assign n30573_o = rb[16];
  assign n30574_o = rb[17];
  assign n30575_o = rb[18];
  assign n30576_o = rb[19];
  assign n30577_o = rb[20];
  /* logical.vhdl:61:45  */
  assign n30578_o = rb[21];
  assign n30579_o = rb[22];
  /* logical.vhdl:61:42  */
  assign n30580_o = rb[23];
  assign n30581_o = rb[24];
  /* logical.vhdl:61:39  */
  assign n30582_o = rb[25];
  assign n30583_o = rb[26];
  /* logical.vhdl:61:36  */
  assign n30584_o = rb[27];
  assign n30585_o = rb[28];
  /* logical.vhdl:61:33  */
  assign n30586_o = rb[29];
  assign n30587_o = rb[30];
  /* logical.vhdl:61:30  */
  assign n30588_o = rb[31];
  assign n30589_o = rb[32];
  /* logical.vhdl:61:27  */
  assign n30590_o = rb[33];
  assign n30591_o = rb[34];
  /* logical.vhdl:61:24  */
  assign n30592_o = rb[35];
  assign n30593_o = rb[36];
  /* logical.vhdl:61:21  */
  assign n30594_o = rb[37];
  assign n30595_o = rb[38];
  /* logical.vhdl:61:18  */
  assign n30596_o = rb[39];
  assign n30597_o = rb[40];
  /* logical.vhdl:60:18  */
  assign n30598_o = rb[41];
  assign n30599_o = rb[42];
  /* logical.vhdl:59:14  */
  assign n30600_o = rb[43];
  /* logical.vhdl:59:14  */
  assign n30601_o = rb[44];
  assign n30602_o = rb[45];
  /* logical.vhdl:59:14  */
  assign n30603_o = rb[46];
  assign n30604_o = rb[47];
  assign n30605_o = rb[48];
  assign n30606_o = rb[49];
  assign n30607_o = rb[50];
  assign n30608_o = rb[51];
  assign n30609_o = rb[52];
  assign n30610_o = rb[53];
  assign n30611_o = rb[54];
  assign n30612_o = rb[55];
  assign n30613_o = rb[56];
  assign n30614_o = rb[57];
  assign n30615_o = rb[58];
  assign n30616_o = rb[59];
  assign n30617_o = rb[60];
  assign n30618_o = rb[61];
  assign n30619_o = rb[62];
  assign n30620_o = rb[63];
  /* logical.vhdl:114:33  */
  assign n30621_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30621_o)
      2'b00: n30622_o = n30557_o;
      2'b01: n30622_o = n30558_o;
      2'b10: n30622_o = n30559_o;
      2'b11: n30622_o = n30560_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30623_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30623_o)
      2'b00: n30624_o = n30561_o;
      2'b01: n30624_o = n30562_o;
      2'b10: n30624_o = n30563_o;
      2'b11: n30624_o = n30564_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30625_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30625_o)
      2'b00: n30626_o = n30565_o;
      2'b01: n30626_o = n30566_o;
      2'b10: n30626_o = n30567_o;
      2'b11: n30626_o = n30568_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30627_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30627_o)
      2'b00: n30628_o = n30569_o;
      2'b01: n30628_o = n30570_o;
      2'b10: n30628_o = n30571_o;
      2'b11: n30628_o = n30572_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30629_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30629_o)
      2'b00: n30630_o = n30573_o;
      2'b01: n30630_o = n30574_o;
      2'b10: n30630_o = n30575_o;
      2'b11: n30630_o = n30576_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30631_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30631_o)
      2'b00: n30632_o = n30577_o;
      2'b01: n30632_o = n30578_o;
      2'b10: n30632_o = n30579_o;
      2'b11: n30632_o = n30580_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30633_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30633_o)
      2'b00: n30634_o = n30581_o;
      2'b01: n30634_o = n30582_o;
      2'b10: n30634_o = n30583_o;
      2'b11: n30634_o = n30584_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30635_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30635_o)
      2'b00: n30636_o = n30585_o;
      2'b01: n30636_o = n30586_o;
      2'b10: n30636_o = n30587_o;
      2'b11: n30636_o = n30588_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30637_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30637_o)
      2'b00: n30638_o = n30589_o;
      2'b01: n30638_o = n30590_o;
      2'b10: n30638_o = n30591_o;
      2'b11: n30638_o = n30592_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30639_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30639_o)
      2'b00: n30640_o = n30593_o;
      2'b01: n30640_o = n30594_o;
      2'b10: n30640_o = n30595_o;
      2'b11: n30640_o = n30596_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30641_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30641_o)
      2'b00: n30642_o = n30597_o;
      2'b01: n30642_o = n30598_o;
      2'b10: n30642_o = n30599_o;
      2'b11: n30642_o = n30600_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30643_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30643_o)
      2'b00: n30644_o = n30601_o;
      2'b01: n30644_o = n30602_o;
      2'b10: n30644_o = n30603_o;
      2'b11: n30644_o = n30604_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30645_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30645_o)
      2'b00: n30646_o = n30605_o;
      2'b01: n30646_o = n30606_o;
      2'b10: n30646_o = n30607_o;
      2'b11: n30646_o = n30608_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30647_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30647_o)
      2'b00: n30648_o = n30609_o;
      2'b01: n30648_o = n30610_o;
      2'b10: n30648_o = n30611_o;
      2'b11: n30648_o = n30612_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30649_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30649_o)
      2'b00: n30650_o = n30613_o;
      2'b01: n30650_o = n30614_o;
      2'b10: n30650_o = n30615_o;
      2'b11: n30650_o = n30616_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30651_o = n28954_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30651_o)
      2'b00: n30652_o = n30617_o;
      2'b01: n30652_o = n30618_o;
      2'b10: n30652_o = n30619_o;
      2'b11: n30652_o = n30620_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30653_o = n28954_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30653_o)
      2'b00: n30654_o = n30622_o;
      2'b01: n30654_o = n30624_o;
      2'b10: n30654_o = n30626_o;
      2'b11: n30654_o = n30628_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30655_o = n28954_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30655_o)
      2'b00: n30656_o = n30630_o;
      2'b01: n30656_o = n30632_o;
      2'b10: n30656_o = n30634_o;
      2'b11: n30656_o = n30636_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30657_o = n28954_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30657_o)
      2'b00: n30658_o = n30638_o;
      2'b01: n30658_o = n30640_o;
      2'b10: n30658_o = n30642_o;
      2'b11: n30658_o = n30644_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30659_o = n28954_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30659_o)
      2'b00: n30660_o = n30646_o;
      2'b01: n30660_o = n30648_o;
      2'b10: n30660_o = n30650_o;
      2'b11: n30660_o = n30652_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30661_o = n28954_o[5:4];
  /* logical.vhdl:114:33  */
  always @*
    case (n30661_o)
      2'b00: n30662_o = n30654_o;
      2'b01: n30662_o = n30656_o;
      2'b10: n30662_o = n30658_o;
      2'b11: n30662_o = n30660_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30663_o = rb[0];
  /* logical.vhdl:114:34  */
  assign n30664_o = rb[1];
  assign n30665_o = rb[2];
  assign n30666_o = rb[3];
  assign n30667_o = rb[4];
  assign n30668_o = rb[5];
  assign n30669_o = rb[6];
  assign n30670_o = rb[7];
  assign n30671_o = rb[8];
  assign n30672_o = rb[9];
  assign n30673_o = rb[10];
  assign n30674_o = rb[11];
  assign n30675_o = rb[12];
  /* logical.vhdl:29:51  */
  assign n30676_o = rb[13];
  assign n30677_o = rb[14];
  /* logical.vhdl:29:48  */
  assign n30678_o = rb[15];
  assign n30679_o = rb[16];
  /* logical.vhdl:29:45  */
  assign n30680_o = rb[17];
  assign n30681_o = rb[18];
  /* logical.vhdl:29:42  */
  assign n30682_o = rb[19];
  assign n30683_o = rb[20];
  /* logical.vhdl:29:39  */
  assign n30684_o = rb[21];
  assign n30685_o = rb[22];
  /* logical.vhdl:29:36  */
  assign n30686_o = rb[23];
  assign n30687_o = rb[24];
  /* logical.vhdl:29:33  */
  assign n30688_o = rb[25];
  assign n30689_o = rb[26];
  /* logical.vhdl:29:30  */
  assign n30690_o = rb[27];
  assign n30691_o = rb[28];
  /* logical.vhdl:29:27  */
  assign n30692_o = rb[29];
  assign n30693_o = rb[30];
  /* logical.vhdl:29:24  */
  assign n30694_o = rb[31];
  assign n30695_o = rb[32];
  /* logical.vhdl:29:21  */
  assign n30696_o = rb[33];
  assign n30697_o = rb[34];
  /* logical.vhdl:29:18  */
  assign n30698_o = rb[35];
  assign n30699_o = rb[36];
  /* logical.vhdl:28:18  */
  assign n30700_o = rb[37];
  assign n30701_o = rb[38];
  /* logical.vhdl:27:14  */
  assign n30702_o = rb[39];
  /* logical.vhdl:27:14  */
  assign n30703_o = rb[40];
  assign n30704_o = rb[41];
  /* logical.vhdl:27:14  */
  assign n30705_o = rb[42];
  assign n30706_o = rb[43];
  assign n30707_o = rb[44];
  assign n30708_o = rb[45];
  assign n30709_o = rb[46];
  assign n30710_o = rb[47];
  assign n30711_o = rb[48];
  assign n30712_o = rb[49];
  assign n30713_o = rb[50];
  assign n30714_o = rb[51];
  assign n30715_o = rb[52];
  assign n30716_o = rb[53];
  assign n30717_o = rb[54];
  assign n30718_o = rb[55];
  assign n30719_o = rb[56];
  assign n30720_o = rb[57];
  assign n30721_o = rb[58];
  assign n30722_o = rb[59];
  assign n30723_o = rb[60];
  assign n30724_o = rb[61];
  assign n30725_o = rb[62];
  assign n30726_o = rb[63];
  /* logical.vhdl:114:33  */
  assign n30727_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30727_o)
      2'b00: n30728_o = n30663_o;
      2'b01: n30728_o = n30664_o;
      2'b10: n30728_o = n30665_o;
      2'b11: n30728_o = n30666_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30729_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30729_o)
      2'b00: n30730_o = n30667_o;
      2'b01: n30730_o = n30668_o;
      2'b10: n30730_o = n30669_o;
      2'b11: n30730_o = n30670_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30731_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30731_o)
      2'b00: n30732_o = n30671_o;
      2'b01: n30732_o = n30672_o;
      2'b10: n30732_o = n30673_o;
      2'b11: n30732_o = n30674_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30733_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30733_o)
      2'b00: n30734_o = n30675_o;
      2'b01: n30734_o = n30676_o;
      2'b10: n30734_o = n30677_o;
      2'b11: n30734_o = n30678_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30735_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30735_o)
      2'b00: n30736_o = n30679_o;
      2'b01: n30736_o = n30680_o;
      2'b10: n30736_o = n30681_o;
      2'b11: n30736_o = n30682_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30737_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30737_o)
      2'b00: n30738_o = n30683_o;
      2'b01: n30738_o = n30684_o;
      2'b10: n30738_o = n30685_o;
      2'b11: n30738_o = n30686_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30739_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30739_o)
      2'b00: n30740_o = n30687_o;
      2'b01: n30740_o = n30688_o;
      2'b10: n30740_o = n30689_o;
      2'b11: n30740_o = n30690_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30741_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30741_o)
      2'b00: n30742_o = n30691_o;
      2'b01: n30742_o = n30692_o;
      2'b10: n30742_o = n30693_o;
      2'b11: n30742_o = n30694_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30743_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30743_o)
      2'b00: n30744_o = n30695_o;
      2'b01: n30744_o = n30696_o;
      2'b10: n30744_o = n30697_o;
      2'b11: n30744_o = n30698_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30745_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30745_o)
      2'b00: n30746_o = n30699_o;
      2'b01: n30746_o = n30700_o;
      2'b10: n30746_o = n30701_o;
      2'b11: n30746_o = n30702_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30747_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30747_o)
      2'b00: n30748_o = n30703_o;
      2'b01: n30748_o = n30704_o;
      2'b10: n30748_o = n30705_o;
      2'b11: n30748_o = n30706_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30749_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30749_o)
      2'b00: n30750_o = n30707_o;
      2'b01: n30750_o = n30708_o;
      2'b10: n30750_o = n30709_o;
      2'b11: n30750_o = n30710_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30751_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30751_o)
      2'b00: n30752_o = n30711_o;
      2'b01: n30752_o = n30712_o;
      2'b10: n30752_o = n30713_o;
      2'b11: n30752_o = n30714_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30753_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30753_o)
      2'b00: n30754_o = n30715_o;
      2'b01: n30754_o = n30716_o;
      2'b10: n30754_o = n30717_o;
      2'b11: n30754_o = n30718_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30755_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30755_o)
      2'b00: n30756_o = n30719_o;
      2'b01: n30756_o = n30720_o;
      2'b10: n30756_o = n30721_o;
      2'b11: n30756_o = n30722_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30757_o = n28964_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30757_o)
      2'b00: n30758_o = n30723_o;
      2'b01: n30758_o = n30724_o;
      2'b10: n30758_o = n30725_o;
      2'b11: n30758_o = n30726_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30759_o = n28964_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30759_o)
      2'b00: n30760_o = n30728_o;
      2'b01: n30760_o = n30730_o;
      2'b10: n30760_o = n30732_o;
      2'b11: n30760_o = n30734_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30761_o = n28964_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30761_o)
      2'b00: n30762_o = n30736_o;
      2'b01: n30762_o = n30738_o;
      2'b10: n30762_o = n30740_o;
      2'b11: n30762_o = n30742_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30763_o = n28964_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30763_o)
      2'b00: n30764_o = n30744_o;
      2'b01: n30764_o = n30746_o;
      2'b10: n30764_o = n30748_o;
      2'b11: n30764_o = n30750_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30765_o = n28964_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30765_o)
      2'b00: n30766_o = n30752_o;
      2'b01: n30766_o = n30754_o;
      2'b10: n30766_o = n30756_o;
      2'b11: n30766_o = n30758_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30767_o = n28964_o[5:4];
  /* logical.vhdl:114:33  */
  always @*
    case (n30767_o)
      2'b00: n30768_o = n30760_o;
      2'b01: n30768_o = n30762_o;
      2'b10: n30768_o = n30764_o;
      2'b11: n30768_o = n30766_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30769_o = rb[0];
  /* logical.vhdl:114:34  */
  assign n30770_o = rb[1];
  assign n30771_o = rb[2];
  assign n30772_o = rb[3];
  assign n30773_o = rb[4];
  assign n30774_o = rb[5];
  assign n30775_o = rb[6];
  assign n30776_o = rb[7];
  assign n30777_o = rb[8];
  assign n30778_o = rb[9];
  assign n30779_o = rb[10];
  assign n30780_o = rb[11];
  assign n30781_o = rb[12];
  /* logical.vhdl:29:51  */
  assign n30782_o = rb[13];
  assign n30783_o = rb[14];
  /* logical.vhdl:29:48  */
  assign n30784_o = rb[15];
  assign n30785_o = rb[16];
  /* logical.vhdl:29:45  */
  assign n30786_o = rb[17];
  assign n30787_o = rb[18];
  /* logical.vhdl:29:42  */
  assign n30788_o = rb[19];
  assign n30789_o = rb[20];
  /* logical.vhdl:29:39  */
  assign n30790_o = rb[21];
  assign n30791_o = rb[22];
  /* logical.vhdl:29:36  */
  assign n30792_o = rb[23];
  assign n30793_o = rb[24];
  /* logical.vhdl:29:33  */
  assign n30794_o = rb[25];
  assign n30795_o = rb[26];
  /* logical.vhdl:29:30  */
  assign n30796_o = rb[27];
  assign n30797_o = rb[28];
  /* logical.vhdl:29:27  */
  assign n30798_o = rb[29];
  assign n30799_o = rb[30];
  /* logical.vhdl:29:24  */
  assign n30800_o = rb[31];
  assign n30801_o = rb[32];
  /* logical.vhdl:29:21  */
  assign n30802_o = rb[33];
  assign n30803_o = rb[34];
  /* logical.vhdl:29:18  */
  assign n30804_o = rb[35];
  assign n30805_o = rb[36];
  /* logical.vhdl:28:18  */
  assign n30806_o = rb[37];
  assign n30807_o = rb[38];
  /* logical.vhdl:27:14  */
  assign n30808_o = rb[39];
  /* logical.vhdl:27:14  */
  assign n30809_o = rb[40];
  assign n30810_o = rb[41];
  /* logical.vhdl:27:14  */
  assign n30811_o = rb[42];
  assign n30812_o = rb[43];
  assign n30813_o = rb[44];
  assign n30814_o = rb[45];
  assign n30815_o = rb[46];
  assign n30816_o = rb[47];
  assign n30817_o = rb[48];
  assign n30818_o = rb[49];
  assign n30819_o = rb[50];
  assign n30820_o = rb[51];
  assign n30821_o = rb[52];
  assign n30822_o = rb[53];
  assign n30823_o = rb[54];
  assign n30824_o = rb[55];
  assign n30825_o = rb[56];
  assign n30826_o = rb[57];
  assign n30827_o = rb[58];
  assign n30828_o = rb[59];
  assign n30829_o = rb[60];
  assign n30830_o = rb[61];
  assign n30831_o = rb[62];
  assign n30832_o = rb[63];
  /* logical.vhdl:114:33  */
  assign n30833_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30833_o)
      2'b00: n30834_o = n30769_o;
      2'b01: n30834_o = n30770_o;
      2'b10: n30834_o = n30771_o;
      2'b11: n30834_o = n30772_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30835_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30835_o)
      2'b00: n30836_o = n30773_o;
      2'b01: n30836_o = n30774_o;
      2'b10: n30836_o = n30775_o;
      2'b11: n30836_o = n30776_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30837_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30837_o)
      2'b00: n30838_o = n30777_o;
      2'b01: n30838_o = n30778_o;
      2'b10: n30838_o = n30779_o;
      2'b11: n30838_o = n30780_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30839_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30839_o)
      2'b00: n30840_o = n30781_o;
      2'b01: n30840_o = n30782_o;
      2'b10: n30840_o = n30783_o;
      2'b11: n30840_o = n30784_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30841_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30841_o)
      2'b00: n30842_o = n30785_o;
      2'b01: n30842_o = n30786_o;
      2'b10: n30842_o = n30787_o;
      2'b11: n30842_o = n30788_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30843_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30843_o)
      2'b00: n30844_o = n30789_o;
      2'b01: n30844_o = n30790_o;
      2'b10: n30844_o = n30791_o;
      2'b11: n30844_o = n30792_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30845_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30845_o)
      2'b00: n30846_o = n30793_o;
      2'b01: n30846_o = n30794_o;
      2'b10: n30846_o = n30795_o;
      2'b11: n30846_o = n30796_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30847_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30847_o)
      2'b00: n30848_o = n30797_o;
      2'b01: n30848_o = n30798_o;
      2'b10: n30848_o = n30799_o;
      2'b11: n30848_o = n30800_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30849_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30849_o)
      2'b00: n30850_o = n30801_o;
      2'b01: n30850_o = n30802_o;
      2'b10: n30850_o = n30803_o;
      2'b11: n30850_o = n30804_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30851_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30851_o)
      2'b00: n30852_o = n30805_o;
      2'b01: n30852_o = n30806_o;
      2'b10: n30852_o = n30807_o;
      2'b11: n30852_o = n30808_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30853_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30853_o)
      2'b00: n30854_o = n30809_o;
      2'b01: n30854_o = n30810_o;
      2'b10: n30854_o = n30811_o;
      2'b11: n30854_o = n30812_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30855_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30855_o)
      2'b00: n30856_o = n30813_o;
      2'b01: n30856_o = n30814_o;
      2'b10: n30856_o = n30815_o;
      2'b11: n30856_o = n30816_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30857_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30857_o)
      2'b00: n30858_o = n30817_o;
      2'b01: n30858_o = n30818_o;
      2'b10: n30858_o = n30819_o;
      2'b11: n30858_o = n30820_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30859_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30859_o)
      2'b00: n30860_o = n30821_o;
      2'b01: n30860_o = n30822_o;
      2'b10: n30860_o = n30823_o;
      2'b11: n30860_o = n30824_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30861_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30861_o)
      2'b00: n30862_o = n30825_o;
      2'b01: n30862_o = n30826_o;
      2'b10: n30862_o = n30827_o;
      2'b11: n30862_o = n30828_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30863_o = n28974_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30863_o)
      2'b00: n30864_o = n30829_o;
      2'b01: n30864_o = n30830_o;
      2'b10: n30864_o = n30831_o;
      2'b11: n30864_o = n30832_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30865_o = n28974_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30865_o)
      2'b00: n30866_o = n30834_o;
      2'b01: n30866_o = n30836_o;
      2'b10: n30866_o = n30838_o;
      2'b11: n30866_o = n30840_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30867_o = n28974_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30867_o)
      2'b00: n30868_o = n30842_o;
      2'b01: n30868_o = n30844_o;
      2'b10: n30868_o = n30846_o;
      2'b11: n30868_o = n30848_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30869_o = n28974_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30869_o)
      2'b00: n30870_o = n30850_o;
      2'b01: n30870_o = n30852_o;
      2'b10: n30870_o = n30854_o;
      2'b11: n30870_o = n30856_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30871_o = n28974_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30871_o)
      2'b00: n30872_o = n30858_o;
      2'b01: n30872_o = n30860_o;
      2'b10: n30872_o = n30862_o;
      2'b11: n30872_o = n30864_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30873_o = n28974_o[5:4];
  /* logical.vhdl:114:33  */
  always @*
    case (n30873_o)
      2'b00: n30874_o = n30866_o;
      2'b01: n30874_o = n30868_o;
      2'b10: n30874_o = n30870_o;
      2'b11: n30874_o = n30872_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30875_o = rb[0];
  /* logical.vhdl:114:34  */
  assign n30876_o = rb[1];
  /* helpers.vhdl:18:14  */
  assign n30877_o = rb[2];
  /* helpers.vhdl:18:14  */
  assign n30878_o = rb[3];
  assign n30879_o = rb[4];
  /* helpers.vhdl:18:14  */
  assign n30880_o = rb[5];
  assign n30881_o = rb[6];
  assign n30882_o = rb[7];
  /* helpers.vhdl:124:18  */
  assign n30883_o = rb[8];
  assign n30884_o = rb[9];
  /* helpers.vhdl:18:14  */
  assign n30885_o = rb[10];
  /* helpers.vhdl:18:14  */
  assign n30886_o = rb[11];
  assign n30887_o = rb[12];
  /* helpers.vhdl:18:14  */
  assign n30888_o = rb[13];
  assign n30889_o = rb[14];
  assign n30890_o = rb[15];
  /* helpers.vhdl:124:18  */
  assign n30891_o = rb[16];
  assign n30892_o = rb[17];
  /* helpers.vhdl:18:14  */
  assign n30893_o = rb[18];
  /* helpers.vhdl:18:14  */
  assign n30894_o = rb[19];
  assign n30895_o = rb[20];
  /* helpers.vhdl:18:14  */
  assign n30896_o = rb[21];
  assign n30897_o = rb[22];
  assign n30898_o = rb[23];
  /* helpers.vhdl:124:18  */
  assign n30899_o = rb[24];
  assign n30900_o = rb[25];
  /* helpers.vhdl:18:14  */
  assign n30901_o = rb[26];
  /* helpers.vhdl:18:14  */
  assign n30902_o = rb[27];
  assign n30903_o = rb[28];
  /* helpers.vhdl:18:14  */
  assign n30904_o = rb[29];
  assign n30905_o = rb[30];
  assign n30906_o = rb[31];
  /* helpers.vhdl:124:18  */
  assign n30907_o = rb[32];
  assign n30908_o = rb[33];
  /* helpers.vhdl:18:14  */
  assign n30909_o = rb[34];
  /* helpers.vhdl:18:14  */
  assign n30910_o = rb[35];
  assign n30911_o = rb[36];
  /* helpers.vhdl:18:14  */
  assign n30912_o = rb[37];
  assign n30913_o = rb[38];
  assign n30914_o = rb[39];
  /* helpers.vhdl:124:18  */
  assign n30915_o = rb[40];
  assign n30916_o = rb[41];
  /* helpers.vhdl:18:14  */
  assign n30917_o = rb[42];
  /* helpers.vhdl:18:14  */
  assign n30918_o = rb[43];
  assign n30919_o = rb[44];
  /* helpers.vhdl:18:14  */
  assign n30920_o = rb[45];
  assign n30921_o = rb[46];
  assign n30922_o = rb[47];
  assign n30923_o = rb[48];
  /* helpers.vhdl:124:18  */
  assign n30924_o = rb[49];
  assign n30925_o = rb[50];
  /* helpers.vhdl:18:14  */
  assign n30926_o = rb[51];
  /* helpers.vhdl:18:14  */
  assign n30927_o = rb[52];
  assign n30928_o = rb[53];
  /* helpers.vhdl:18:14  */
  assign n30929_o = rb[54];
  /* ppc_fx_insns.vhdl:740:26  */
  assign n30930_o = rb[55];
  assign n30931_o = rb[56];
  /* ppc_fx_insns.vhdl:739:26  */
  assign n30932_o = rb[57];
  assign n30933_o = rb[58];
  /* ppc_fx_insns.vhdl:738:26  */
  assign n30934_o = rb[59];
  assign n30935_o = rb[60];
  /* ppc_fx_insns.vhdl:89:18  */
  assign n30936_o = rb[61];
  /* ppc_fx_insns.vhdl:89:18  */
  assign n30937_o = rb[62];
  assign n30938_o = rb[63];
  /* logical.vhdl:114:33  */
  assign n30939_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30939_o)
      2'b00: n30940_o = n30875_o;
      2'b01: n30940_o = n30876_o;
      2'b10: n30940_o = n30877_o;
      2'b11: n30940_o = n30878_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30941_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30941_o)
      2'b00: n30942_o = n30879_o;
      2'b01: n30942_o = n30880_o;
      2'b10: n30942_o = n30881_o;
      2'b11: n30942_o = n30882_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30943_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30943_o)
      2'b00: n30944_o = n30883_o;
      2'b01: n30944_o = n30884_o;
      2'b10: n30944_o = n30885_o;
      2'b11: n30944_o = n30886_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30945_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30945_o)
      2'b00: n30946_o = n30887_o;
      2'b01: n30946_o = n30888_o;
      2'b10: n30946_o = n30889_o;
      2'b11: n30946_o = n30890_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30947_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30947_o)
      2'b00: n30948_o = n30891_o;
      2'b01: n30948_o = n30892_o;
      2'b10: n30948_o = n30893_o;
      2'b11: n30948_o = n30894_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30949_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30949_o)
      2'b00: n30950_o = n30895_o;
      2'b01: n30950_o = n30896_o;
      2'b10: n30950_o = n30897_o;
      2'b11: n30950_o = n30898_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30951_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30951_o)
      2'b00: n30952_o = n30899_o;
      2'b01: n30952_o = n30900_o;
      2'b10: n30952_o = n30901_o;
      2'b11: n30952_o = n30902_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30953_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30953_o)
      2'b00: n30954_o = n30903_o;
      2'b01: n30954_o = n30904_o;
      2'b10: n30954_o = n30905_o;
      2'b11: n30954_o = n30906_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30955_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30955_o)
      2'b00: n30956_o = n30907_o;
      2'b01: n30956_o = n30908_o;
      2'b10: n30956_o = n30909_o;
      2'b11: n30956_o = n30910_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30957_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30957_o)
      2'b00: n30958_o = n30911_o;
      2'b01: n30958_o = n30912_o;
      2'b10: n30958_o = n30913_o;
      2'b11: n30958_o = n30914_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30959_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30959_o)
      2'b00: n30960_o = n30915_o;
      2'b01: n30960_o = n30916_o;
      2'b10: n30960_o = n30917_o;
      2'b11: n30960_o = n30918_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30961_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30961_o)
      2'b00: n30962_o = n30919_o;
      2'b01: n30962_o = n30920_o;
      2'b10: n30962_o = n30921_o;
      2'b11: n30962_o = n30922_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30963_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30963_o)
      2'b00: n30964_o = n30923_o;
      2'b01: n30964_o = n30924_o;
      2'b10: n30964_o = n30925_o;
      2'b11: n30964_o = n30926_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30965_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30965_o)
      2'b00: n30966_o = n30927_o;
      2'b01: n30966_o = n30928_o;
      2'b10: n30966_o = n30929_o;
      2'b11: n30966_o = n30930_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30967_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30967_o)
      2'b00: n30968_o = n30931_o;
      2'b01: n30968_o = n30932_o;
      2'b10: n30968_o = n30933_o;
      2'b11: n30968_o = n30934_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30969_o = n28984_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n30969_o)
      2'b00: n30970_o = n30935_o;
      2'b01: n30970_o = n30936_o;
      2'b10: n30970_o = n30937_o;
      2'b11: n30970_o = n30938_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30971_o = n28984_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30971_o)
      2'b00: n30972_o = n30940_o;
      2'b01: n30972_o = n30942_o;
      2'b10: n30972_o = n30944_o;
      2'b11: n30972_o = n30946_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30973_o = n28984_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30973_o)
      2'b00: n30974_o = n30948_o;
      2'b01: n30974_o = n30950_o;
      2'b10: n30974_o = n30952_o;
      2'b11: n30974_o = n30954_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30975_o = n28984_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30975_o)
      2'b00: n30976_o = n30956_o;
      2'b01: n30976_o = n30958_o;
      2'b10: n30976_o = n30960_o;
      2'b11: n30976_o = n30962_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30977_o = n28984_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n30977_o)
      2'b00: n30978_o = n30964_o;
      2'b01: n30978_o = n30966_o;
      2'b10: n30978_o = n30968_o;
      2'b11: n30978_o = n30970_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30979_o = n28984_o[5:4];
  /* logical.vhdl:114:33  */
  always @*
    case (n30979_o)
      2'b00: n30980_o = n30972_o;
      2'b01: n30980_o = n30974_o;
      2'b10: n30980_o = n30976_o;
      2'b11: n30980_o = n30978_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n30981_o = rb[0];
  /* logical.vhdl:114:34  */
  assign n30982_o = rb[1];
  assign n30983_o = rb[2];
  assign n30984_o = rb[3];
  assign n30985_o = rb[4];
  assign n30986_o = rb[5];
  assign n30987_o = rb[6];
  assign n30988_o = rb[7];
  assign n30989_o = rb[8];
  assign n30990_o = rb[9];
  assign n30991_o = rb[10];
  assign n30992_o = rb[11];
  assign n30993_o = rb[12];
  assign n30994_o = rb[13];
  assign n30995_o = rb[14];
  assign n30996_o = rb[15];
  assign n30997_o = rb[16];
  assign n30998_o = rb[17];
  assign n30999_o = rb[18];
  assign n31000_o = rb[19];
  assign n31001_o = rb[20];
  assign n31002_o = rb[21];
  assign n31003_o = rb[22];
  assign n31004_o = rb[23];
  assign n31005_o = rb[24];
  assign n31006_o = rb[25];
  assign n31007_o = rb[26];
  assign n31008_o = rb[27];
  assign n31009_o = rb[28];
  assign n31010_o = rb[29];
  assign n31011_o = rb[30];
  assign n31012_o = rb[31];
  assign n31013_o = rb[32];
  assign n31014_o = rb[33];
  assign n31015_o = rb[34];
  assign n31016_o = rb[35];
  assign n31017_o = rb[36];
  assign n31018_o = rb[37];
  assign n31019_o = rb[38];
  assign n31020_o = rb[39];
  assign n31021_o = rb[40];
  assign n31022_o = rb[41];
  assign n31023_o = rb[42];
  assign n31024_o = rb[43];
  assign n31025_o = rb[44];
  assign n31026_o = rb[45];
  assign n31027_o = rb[46];
  assign n31028_o = rb[47];
  assign n31029_o = rb[48];
  assign n31030_o = rb[49];
  assign n31031_o = rb[50];
  assign n31032_o = rb[51];
  assign n31033_o = rb[52];
  assign n31034_o = rb[53];
  assign n31035_o = rb[54];
  assign n31036_o = rb[55];
  assign n31037_o = rb[56];
  assign n31038_o = rb[57];
  assign n31039_o = rb[58];
  assign n31040_o = rb[59];
  assign n31041_o = rb[60];
  assign n31042_o = rb[61];
  assign n31043_o = rb[62];
  assign n31044_o = rb[63];
  /* logical.vhdl:114:33  */
  assign n31045_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31045_o)
      2'b00: n31046_o = n30981_o;
      2'b01: n31046_o = n30982_o;
      2'b10: n31046_o = n30983_o;
      2'b11: n31046_o = n30984_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31047_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31047_o)
      2'b00: n31048_o = n30985_o;
      2'b01: n31048_o = n30986_o;
      2'b10: n31048_o = n30987_o;
      2'b11: n31048_o = n30988_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31049_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31049_o)
      2'b00: n31050_o = n30989_o;
      2'b01: n31050_o = n30990_o;
      2'b10: n31050_o = n30991_o;
      2'b11: n31050_o = n30992_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31051_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31051_o)
      2'b00: n31052_o = n30993_o;
      2'b01: n31052_o = n30994_o;
      2'b10: n31052_o = n30995_o;
      2'b11: n31052_o = n30996_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31053_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31053_o)
      2'b00: n31054_o = n30997_o;
      2'b01: n31054_o = n30998_o;
      2'b10: n31054_o = n30999_o;
      2'b11: n31054_o = n31000_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31055_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31055_o)
      2'b00: n31056_o = n31001_o;
      2'b01: n31056_o = n31002_o;
      2'b10: n31056_o = n31003_o;
      2'b11: n31056_o = n31004_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31057_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31057_o)
      2'b00: n31058_o = n31005_o;
      2'b01: n31058_o = n31006_o;
      2'b10: n31058_o = n31007_o;
      2'b11: n31058_o = n31008_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31059_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31059_o)
      2'b00: n31060_o = n31009_o;
      2'b01: n31060_o = n31010_o;
      2'b10: n31060_o = n31011_o;
      2'b11: n31060_o = n31012_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31061_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31061_o)
      2'b00: n31062_o = n31013_o;
      2'b01: n31062_o = n31014_o;
      2'b10: n31062_o = n31015_o;
      2'b11: n31062_o = n31016_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31063_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31063_o)
      2'b00: n31064_o = n31017_o;
      2'b01: n31064_o = n31018_o;
      2'b10: n31064_o = n31019_o;
      2'b11: n31064_o = n31020_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31065_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31065_o)
      2'b00: n31066_o = n31021_o;
      2'b01: n31066_o = n31022_o;
      2'b10: n31066_o = n31023_o;
      2'b11: n31066_o = n31024_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31067_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31067_o)
      2'b00: n31068_o = n31025_o;
      2'b01: n31068_o = n31026_o;
      2'b10: n31068_o = n31027_o;
      2'b11: n31068_o = n31028_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31069_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31069_o)
      2'b00: n31070_o = n31029_o;
      2'b01: n31070_o = n31030_o;
      2'b10: n31070_o = n31031_o;
      2'b11: n31070_o = n31032_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31071_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31071_o)
      2'b00: n31072_o = n31033_o;
      2'b01: n31072_o = n31034_o;
      2'b10: n31072_o = n31035_o;
      2'b11: n31072_o = n31036_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31073_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31073_o)
      2'b00: n31074_o = n31037_o;
      2'b01: n31074_o = n31038_o;
      2'b10: n31074_o = n31039_o;
      2'b11: n31074_o = n31040_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31075_o = n28994_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31075_o)
      2'b00: n31076_o = n31041_o;
      2'b01: n31076_o = n31042_o;
      2'b10: n31076_o = n31043_o;
      2'b11: n31076_o = n31044_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31077_o = n28994_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31077_o)
      2'b00: n31078_o = n31046_o;
      2'b01: n31078_o = n31048_o;
      2'b10: n31078_o = n31050_o;
      2'b11: n31078_o = n31052_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31079_o = n28994_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31079_o)
      2'b00: n31080_o = n31054_o;
      2'b01: n31080_o = n31056_o;
      2'b10: n31080_o = n31058_o;
      2'b11: n31080_o = n31060_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31081_o = n28994_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31081_o)
      2'b00: n31082_o = n31062_o;
      2'b01: n31082_o = n31064_o;
      2'b10: n31082_o = n31066_o;
      2'b11: n31082_o = n31068_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31083_o = n28994_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31083_o)
      2'b00: n31084_o = n31070_o;
      2'b01: n31084_o = n31072_o;
      2'b10: n31084_o = n31074_o;
      2'b11: n31084_o = n31076_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31085_o = n28994_o[5:4];
  /* logical.vhdl:114:33  */
  always @*
    case (n31085_o)
      2'b00: n31086_o = n31078_o;
      2'b01: n31086_o = n31080_o;
      2'b10: n31086_o = n31082_o;
      2'b11: n31086_o = n31084_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31087_o = rb[0];
  /* logical.vhdl:114:34  */
  assign n31088_o = rb[1];
  assign n31089_o = rb[2];
  assign n31090_o = rb[3];
  assign n31091_o = rb[4];
  assign n31092_o = rb[5];
  assign n31093_o = rb[6];
  assign n31094_o = rb[7];
  assign n31095_o = rb[8];
  assign n31096_o = rb[9];
  assign n31097_o = rb[10];
  assign n31098_o = rb[11];
  assign n31099_o = rb[12];
  assign n31100_o = rb[13];
  assign n31101_o = rb[14];
  assign n31102_o = rb[15];
  assign n31103_o = rb[16];
  assign n31104_o = rb[17];
  assign n31105_o = rb[18];
  assign n31106_o = rb[19];
  assign n31107_o = rb[20];
  assign n31108_o = rb[21];
  assign n31109_o = rb[22];
  assign n31110_o = rb[23];
  assign n31111_o = rb[24];
  assign n31112_o = rb[25];
  assign n31113_o = rb[26];
  assign n31114_o = rb[27];
  assign n31115_o = rb[28];
  assign n31116_o = rb[29];
  assign n31117_o = rb[30];
  assign n31118_o = rb[31];
  assign n31119_o = rb[32];
  assign n31120_o = rb[33];
  assign n31121_o = rb[34];
  assign n31122_o = rb[35];
  assign n31123_o = rb[36];
  assign n31124_o = rb[37];
  assign n31125_o = rb[38];
  assign n31126_o = rb[39];
  assign n31127_o = rb[40];
  assign n31128_o = rb[41];
  assign n31129_o = rb[42];
  assign n31130_o = rb[43];
  assign n31131_o = rb[44];
  assign n31132_o = rb[45];
  assign n31133_o = rb[46];
  assign n31134_o = rb[47];
  assign n31135_o = rb[48];
  assign n31136_o = rb[49];
  assign n31137_o = rb[50];
  assign n31138_o = rb[51];
  assign n31139_o = rb[52];
  assign n31140_o = rb[53];
  assign n31141_o = rb[54];
  assign n31142_o = rb[55];
  assign n31143_o = rb[56];
  assign n31144_o = rb[57];
  assign n31145_o = rb[58];
  assign n31146_o = rb[59];
  assign n31147_o = rb[60];
  assign n31148_o = rb[61];
  assign n31149_o = rb[62];
  assign n31150_o = rb[63];
  /* logical.vhdl:114:33  */
  assign n31151_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31151_o)
      2'b00: n31152_o = n31087_o;
      2'b01: n31152_o = n31088_o;
      2'b10: n31152_o = n31089_o;
      2'b11: n31152_o = n31090_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31153_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31153_o)
      2'b00: n31154_o = n31091_o;
      2'b01: n31154_o = n31092_o;
      2'b10: n31154_o = n31093_o;
      2'b11: n31154_o = n31094_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31155_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31155_o)
      2'b00: n31156_o = n31095_o;
      2'b01: n31156_o = n31096_o;
      2'b10: n31156_o = n31097_o;
      2'b11: n31156_o = n31098_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31157_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31157_o)
      2'b00: n31158_o = n31099_o;
      2'b01: n31158_o = n31100_o;
      2'b10: n31158_o = n31101_o;
      2'b11: n31158_o = n31102_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31159_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31159_o)
      2'b00: n31160_o = n31103_o;
      2'b01: n31160_o = n31104_o;
      2'b10: n31160_o = n31105_o;
      2'b11: n31160_o = n31106_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31161_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31161_o)
      2'b00: n31162_o = n31107_o;
      2'b01: n31162_o = n31108_o;
      2'b10: n31162_o = n31109_o;
      2'b11: n31162_o = n31110_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31163_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31163_o)
      2'b00: n31164_o = n31111_o;
      2'b01: n31164_o = n31112_o;
      2'b10: n31164_o = n31113_o;
      2'b11: n31164_o = n31114_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31165_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31165_o)
      2'b00: n31166_o = n31115_o;
      2'b01: n31166_o = n31116_o;
      2'b10: n31166_o = n31117_o;
      2'b11: n31166_o = n31118_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31167_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31167_o)
      2'b00: n31168_o = n31119_o;
      2'b01: n31168_o = n31120_o;
      2'b10: n31168_o = n31121_o;
      2'b11: n31168_o = n31122_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31169_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31169_o)
      2'b00: n31170_o = n31123_o;
      2'b01: n31170_o = n31124_o;
      2'b10: n31170_o = n31125_o;
      2'b11: n31170_o = n31126_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31171_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31171_o)
      2'b00: n31172_o = n31127_o;
      2'b01: n31172_o = n31128_o;
      2'b10: n31172_o = n31129_o;
      2'b11: n31172_o = n31130_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31173_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31173_o)
      2'b00: n31174_o = n31131_o;
      2'b01: n31174_o = n31132_o;
      2'b10: n31174_o = n31133_o;
      2'b11: n31174_o = n31134_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31175_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31175_o)
      2'b00: n31176_o = n31135_o;
      2'b01: n31176_o = n31136_o;
      2'b10: n31176_o = n31137_o;
      2'b11: n31176_o = n31138_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31177_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31177_o)
      2'b00: n31178_o = n31139_o;
      2'b01: n31178_o = n31140_o;
      2'b10: n31178_o = n31141_o;
      2'b11: n31178_o = n31142_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31179_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31179_o)
      2'b00: n31180_o = n31143_o;
      2'b01: n31180_o = n31144_o;
      2'b10: n31180_o = n31145_o;
      2'b11: n31180_o = n31146_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31181_o = n29004_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31181_o)
      2'b00: n31182_o = n31147_o;
      2'b01: n31182_o = n31148_o;
      2'b10: n31182_o = n31149_o;
      2'b11: n31182_o = n31150_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31183_o = n29004_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31183_o)
      2'b00: n31184_o = n31152_o;
      2'b01: n31184_o = n31154_o;
      2'b10: n31184_o = n31156_o;
      2'b11: n31184_o = n31158_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31185_o = n29004_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31185_o)
      2'b00: n31186_o = n31160_o;
      2'b01: n31186_o = n31162_o;
      2'b10: n31186_o = n31164_o;
      2'b11: n31186_o = n31166_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31187_o = n29004_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31187_o)
      2'b00: n31188_o = n31168_o;
      2'b01: n31188_o = n31170_o;
      2'b10: n31188_o = n31172_o;
      2'b11: n31188_o = n31174_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31189_o = n29004_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31189_o)
      2'b00: n31190_o = n31176_o;
      2'b01: n31190_o = n31178_o;
      2'b10: n31190_o = n31180_o;
      2'b11: n31190_o = n31182_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31191_o = n29004_o[5:4];
  /* logical.vhdl:114:33  */
  always @*
    case (n31191_o)
      2'b00: n31192_o = n31184_o;
      2'b01: n31192_o = n31186_o;
      2'b10: n31192_o = n31188_o;
      2'b11: n31192_o = n31190_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31193_o = rb[0];
  /* logical.vhdl:114:34  */
  assign n31194_o = rb[1];
  assign n31195_o = rb[2];
  assign n31196_o = rb[3];
  assign n31197_o = rb[4];
  assign n31198_o = rb[5];
  assign n31199_o = rb[6];
  assign n31200_o = rb[7];
  assign n31201_o = rb[8];
  assign n31202_o = rb[9];
  assign n31203_o = rb[10];
  assign n31204_o = rb[11];
  assign n31205_o = rb[12];
  assign n31206_o = rb[13];
  assign n31207_o = rb[14];
  assign n31208_o = rb[15];
  assign n31209_o = rb[16];
  assign n31210_o = rb[17];
  assign n31211_o = rb[18];
  assign n31212_o = rb[19];
  assign n31213_o = rb[20];
  assign n31214_o = rb[21];
  assign n31215_o = rb[22];
  assign n31216_o = rb[23];
  assign n31217_o = rb[24];
  assign n31218_o = rb[25];
  assign n31219_o = rb[26];
  assign n31220_o = rb[27];
  assign n31221_o = rb[28];
  assign n31222_o = rb[29];
  assign n31223_o = rb[30];
  assign n31224_o = rb[31];
  assign n31225_o = rb[32];
  assign n31226_o = rb[33];
  assign n31227_o = rb[34];
  assign n31228_o = rb[35];
  assign n31229_o = rb[36];
  assign n31230_o = rb[37];
  assign n31231_o = rb[38];
  assign n31232_o = rb[39];
  assign n31233_o = rb[40];
  assign n31234_o = rb[41];
  assign n31235_o = rb[42];
  assign n31236_o = rb[43];
  assign n31237_o = rb[44];
  assign n31238_o = rb[45];
  assign n31239_o = rb[46];
  assign n31240_o = rb[47];
  assign n31241_o = rb[48];
  assign n31242_o = rb[49];
  assign n31243_o = rb[50];
  assign n31244_o = rb[51];
  assign n31245_o = rb[52];
  assign n31246_o = rb[53];
  assign n31247_o = rb[54];
  assign n31248_o = rb[55];
  assign n31249_o = rb[56];
  assign n31250_o = rb[57];
  assign n31251_o = rb[58];
  assign n31252_o = rb[59];
  assign n31253_o = rb[60];
  assign n31254_o = rb[61];
  assign n31255_o = rb[62];
  assign n31256_o = rb[63];
  /* logical.vhdl:114:33  */
  assign n31257_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31257_o)
      2'b00: n31258_o = n31193_o;
      2'b01: n31258_o = n31194_o;
      2'b10: n31258_o = n31195_o;
      2'b11: n31258_o = n31196_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31259_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31259_o)
      2'b00: n31260_o = n31197_o;
      2'b01: n31260_o = n31198_o;
      2'b10: n31260_o = n31199_o;
      2'b11: n31260_o = n31200_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31261_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31261_o)
      2'b00: n31262_o = n31201_o;
      2'b01: n31262_o = n31202_o;
      2'b10: n31262_o = n31203_o;
      2'b11: n31262_o = n31204_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31263_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31263_o)
      2'b00: n31264_o = n31205_o;
      2'b01: n31264_o = n31206_o;
      2'b10: n31264_o = n31207_o;
      2'b11: n31264_o = n31208_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31265_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31265_o)
      2'b00: n31266_o = n31209_o;
      2'b01: n31266_o = n31210_o;
      2'b10: n31266_o = n31211_o;
      2'b11: n31266_o = n31212_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31267_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31267_o)
      2'b00: n31268_o = n31213_o;
      2'b01: n31268_o = n31214_o;
      2'b10: n31268_o = n31215_o;
      2'b11: n31268_o = n31216_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31269_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31269_o)
      2'b00: n31270_o = n31217_o;
      2'b01: n31270_o = n31218_o;
      2'b10: n31270_o = n31219_o;
      2'b11: n31270_o = n31220_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31271_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31271_o)
      2'b00: n31272_o = n31221_o;
      2'b01: n31272_o = n31222_o;
      2'b10: n31272_o = n31223_o;
      2'b11: n31272_o = n31224_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31273_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31273_o)
      2'b00: n31274_o = n31225_o;
      2'b01: n31274_o = n31226_o;
      2'b10: n31274_o = n31227_o;
      2'b11: n31274_o = n31228_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31275_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31275_o)
      2'b00: n31276_o = n31229_o;
      2'b01: n31276_o = n31230_o;
      2'b10: n31276_o = n31231_o;
      2'b11: n31276_o = n31232_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31277_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31277_o)
      2'b00: n31278_o = n31233_o;
      2'b01: n31278_o = n31234_o;
      2'b10: n31278_o = n31235_o;
      2'b11: n31278_o = n31236_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31279_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31279_o)
      2'b00: n31280_o = n31237_o;
      2'b01: n31280_o = n31238_o;
      2'b10: n31280_o = n31239_o;
      2'b11: n31280_o = n31240_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31281_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31281_o)
      2'b00: n31282_o = n31241_o;
      2'b01: n31282_o = n31242_o;
      2'b10: n31282_o = n31243_o;
      2'b11: n31282_o = n31244_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31283_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31283_o)
      2'b00: n31284_o = n31245_o;
      2'b01: n31284_o = n31246_o;
      2'b10: n31284_o = n31247_o;
      2'b11: n31284_o = n31248_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31285_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31285_o)
      2'b00: n31286_o = n31249_o;
      2'b01: n31286_o = n31250_o;
      2'b10: n31286_o = n31251_o;
      2'b11: n31286_o = n31252_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31287_o = n29014_o[1:0];
  /* logical.vhdl:114:33  */
  always @*
    case (n31287_o)
      2'b00: n31288_o = n31253_o;
      2'b01: n31288_o = n31254_o;
      2'b10: n31288_o = n31255_o;
      2'b11: n31288_o = n31256_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31289_o = n29014_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31289_o)
      2'b00: n31290_o = n31258_o;
      2'b01: n31290_o = n31260_o;
      2'b10: n31290_o = n31262_o;
      2'b11: n31290_o = n31264_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31291_o = n29014_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31291_o)
      2'b00: n31292_o = n31266_o;
      2'b01: n31292_o = n31268_o;
      2'b10: n31292_o = n31270_o;
      2'b11: n31292_o = n31272_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31293_o = n29014_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31293_o)
      2'b00: n31294_o = n31274_o;
      2'b01: n31294_o = n31276_o;
      2'b10: n31294_o = n31278_o;
      2'b11: n31294_o = n31280_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31295_o = n29014_o[3:2];
  /* logical.vhdl:114:33  */
  always @*
    case (n31295_o)
      2'b00: n31296_o = n31282_o;
      2'b01: n31296_o = n31284_o;
      2'b10: n31296_o = n31286_o;
      2'b11: n31296_o = n31288_o;
    endcase
  /* logical.vhdl:114:33  */
  assign n31297_o = n29014_o[5:4];
  /* logical.vhdl:114:33  */
  always @*
    case (n31297_o)
      2'b00: n31298_o = n31290_o;
      2'b01: n31298_o = n31292_o;
      2'b10: n31298_o = n31294_o;
      2'b11: n31298_o = n31296_o;
    endcase
endmodule

module rotator
  (input  [63:0] rs,
   input  [63:0] ra,
   input  [6:0] shift,
   input  [31:0] insn,
   input  is_32bit,
   input  right_shift,
   input  arith,
   input  clear_left,
   input  clear_right,
   input  sign_ext_rs,
   output [63:0] result,
   output carry_out);
  wire [63:0] repl32;
  wire [5:0] rot_count;
  wire [63:0] rot1;
  wire [63:0] rot2;
  wire [63:0] rot;
  wire [6:0] sh;
  wire [6:0] mb;
  wire [6:0] me;
  wire [63:0] mr;
  wire [63:0] ml;
  wire [1:0] output_mode;
  wire [31:0] n27734_o;
  wire n27735_o;
  wire n27736_o;
  wire n27737_o;
  wire n27738_o;
  wire n27739_o;
  wire n27740_o;
  wire n27741_o;
  wire n27742_o;
  wire n27743_o;
  wire n27744_o;
  wire n27745_o;
  wire n27746_o;
  wire n27747_o;
  wire n27748_o;
  wire n27749_o;
  wire n27750_o;
  wire n27751_o;
  wire n27752_o;
  wire n27753_o;
  wire n27754_o;
  wire n27755_o;
  wire n27756_o;
  wire n27757_o;
  wire n27758_o;
  wire n27759_o;
  wire n27760_o;
  wire n27761_o;
  wire n27762_o;
  wire n27763_o;
  wire n27764_o;
  wire n27765_o;
  wire n27766_o;
  wire [3:0] n27767_o;
  wire [3:0] n27768_o;
  wire [3:0] n27769_o;
  wire [3:0] n27770_o;
  wire [3:0] n27771_o;
  wire [3:0] n27772_o;
  wire [3:0] n27773_o;
  wire [3:0] n27774_o;
  wire [15:0] n27775_o;
  wire [15:0] n27776_o;
  wire [31:0] n27777_o;
  wire [31:0] n27778_o;
  wire [31:0] n27779_o;
  wire [31:0] n27780_o;
  wire [31:0] n27781_o;
  wire [63:0] n27782_o;
  wire [5:0] n27783_o;
  wire [5:0] n27784_o;
  wire [5:0] n27785_o;
  wire [5:0] n27786_o;
  wire [1:0] n27787_o;
  wire n27789_o;
  wire [62:0] n27790_o;
  wire n27791_o;
  wire [63:0] n27792_o;
  wire n27794_o;
  wire [61:0] n27795_o;
  wire [1:0] n27796_o;
  wire [63:0] n27797_o;
  wire n27799_o;
  wire [60:0] n27800_o;
  wire [2:0] n27801_o;
  wire [63:0] n27802_o;
  wire [2:0] n27803_o;
  reg [63:0] n27804_o;
  wire [1:0] n27805_o;
  wire n27807_o;
  wire [59:0] n27808_o;
  wire [3:0] n27809_o;
  wire [63:0] n27810_o;
  wire n27812_o;
  wire [55:0] n27813_o;
  wire [7:0] n27814_o;
  wire [63:0] n27815_o;
  wire n27817_o;
  wire [51:0] n27818_o;
  wire [11:0] n27819_o;
  wire [63:0] n27820_o;
  wire [2:0] n27821_o;
  reg [63:0] n27822_o;
  wire [1:0] n27823_o;
  wire n27825_o;
  wire [47:0] n27826_o;
  wire [15:0] n27827_o;
  wire [63:0] n27828_o;
  wire n27830_o;
  wire [31:0] n27831_o;
  wire [31:0] n27832_o;
  wire [63:0] n27833_o;
  wire n27835_o;
  wire [15:0] n27836_o;
  wire [47:0] n27837_o;
  wire [63:0] n27838_o;
  wire [2:0] n27839_o;
  reg [63:0] n27840_o;
  wire n27841_o;
  wire n27842_o;
  wire n27843_o;
  wire [5:0] n27844_o;
  wire [6:0] n27845_o;
  wire [4:0] n27846_o;
  wire [6:0] n27848_o;
  wire n27849_o;
  wire [1:0] n27851_o;
  wire [4:0] n27852_o;
  wire [6:0] n27853_o;
  wire [6:0] n27854_o;
  wire n27855_o;
  wire n27856_o;
  wire n27857_o;
  wire [1:0] n27858_o;
  wire [4:0] n27859_o;
  wire [6:0] n27860_o;
  wire [6:0] n27861_o;
  wire [1:0] n27863_o;
  wire [6:0] n27865_o;
  wire [6:0] n27866_o;
  wire [6:0] n27867_o;
  wire n27868_o;
  wire [4:0] n27869_o;
  wire [6:0] n27871_o;
  wire n27872_o;
  wire n27873_o;
  wire n27874_o;
  wire [1:0] n27876_o;
  wire [4:0] n27877_o;
  wire [6:0] n27878_o;
  wire n27879_o;
  wire [5:0] n27880_o;
  wire [5:0] n27881_o;
  wire [6:0] n27882_o;
  wire [6:0] n27883_o;
  wire [6:0] n27884_o;
  wire [30:0] n27891_o;
  wire [31:0] n27892_o;
  wire n27894_o;
  wire n27897_o;
  localparam [63:0] n27898_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire [30:0] n27900_o;
  wire [31:0] n27901_o;
  wire n27903_o;
  wire n27905_o;
  wire n27906_o;
  wire [30:0] n27908_o;
  wire [31:0] n27909_o;
  wire n27911_o;
  wire n27913_o;
  wire n27914_o;
  wire [30:0] n27916_o;
  wire [31:0] n27917_o;
  wire n27919_o;
  wire n27921_o;
  wire n27922_o;
  wire [30:0] n27924_o;
  wire [31:0] n27925_o;
  wire n27927_o;
  wire n27929_o;
  wire n27930_o;
  wire [30:0] n27932_o;
  wire [31:0] n27933_o;
  wire n27935_o;
  wire n27937_o;
  wire n27938_o;
  wire [30:0] n27940_o;
  wire [31:0] n27941_o;
  wire n27943_o;
  wire n27945_o;
  wire n27946_o;
  wire [30:0] n27948_o;
  wire [31:0] n27949_o;
  wire n27951_o;
  wire n27953_o;
  wire n27954_o;
  wire [30:0] n27956_o;
  wire [31:0] n27957_o;
  wire n27959_o;
  wire n27961_o;
  wire n27962_o;
  wire [30:0] n27964_o;
  wire [31:0] n27965_o;
  wire n27967_o;
  wire n27969_o;
  wire n27970_o;
  wire [30:0] n27972_o;
  wire [31:0] n27973_o;
  wire n27975_o;
  wire n27977_o;
  wire n27978_o;
  wire [30:0] n27980_o;
  wire [31:0] n27981_o;
  wire n27983_o;
  wire n27985_o;
  wire n27986_o;
  wire [30:0] n27988_o;
  wire [31:0] n27989_o;
  wire n27991_o;
  wire n27993_o;
  wire n27994_o;
  wire [30:0] n27996_o;
  wire [31:0] n27997_o;
  wire n27999_o;
  wire n28001_o;
  wire n28002_o;
  wire [30:0] n28004_o;
  wire [31:0] n28005_o;
  wire n28007_o;
  wire n28009_o;
  wire n28010_o;
  wire [30:0] n28012_o;
  wire [31:0] n28013_o;
  wire n28015_o;
  wire n28017_o;
  wire n28018_o;
  wire [30:0] n28020_o;
  wire [31:0] n28021_o;
  wire n28023_o;
  wire n28025_o;
  wire n28026_o;
  wire [30:0] n28028_o;
  wire [31:0] n28029_o;
  wire n28031_o;
  wire n28033_o;
  wire n28034_o;
  wire [30:0] n28036_o;
  wire [31:0] n28037_o;
  wire n28039_o;
  wire n28041_o;
  wire n28042_o;
  wire [30:0] n28044_o;
  wire [31:0] n28045_o;
  wire n28047_o;
  wire n28049_o;
  wire n28050_o;
  wire [30:0] n28052_o;
  wire [31:0] n28053_o;
  wire n28055_o;
  wire n28057_o;
  wire n28058_o;
  wire [30:0] n28060_o;
  wire [31:0] n28061_o;
  wire n28063_o;
  wire n28065_o;
  wire n28066_o;
  wire [30:0] n28068_o;
  wire [31:0] n28069_o;
  wire n28071_o;
  wire n28073_o;
  wire n28074_o;
  wire [30:0] n28076_o;
  wire [31:0] n28077_o;
  wire n28079_o;
  wire n28081_o;
  wire n28082_o;
  wire [30:0] n28084_o;
  wire [31:0] n28085_o;
  wire n28087_o;
  wire n28089_o;
  wire n28090_o;
  wire [30:0] n28092_o;
  wire [31:0] n28093_o;
  wire n28095_o;
  wire n28097_o;
  wire n28098_o;
  wire [30:0] n28100_o;
  wire [31:0] n28101_o;
  wire n28103_o;
  wire n28105_o;
  wire n28106_o;
  wire [30:0] n28108_o;
  wire [31:0] n28109_o;
  wire n28111_o;
  wire n28113_o;
  wire n28114_o;
  wire [30:0] n28116_o;
  wire [31:0] n28117_o;
  wire n28119_o;
  wire n28121_o;
  wire n28122_o;
  wire [30:0] n28124_o;
  wire [31:0] n28125_o;
  wire n28127_o;
  wire n28129_o;
  wire n28130_o;
  wire [30:0] n28132_o;
  wire [31:0] n28133_o;
  wire n28135_o;
  wire n28137_o;
  wire n28138_o;
  wire [30:0] n28140_o;
  wire [31:0] n28141_o;
  wire n28143_o;
  wire n28145_o;
  wire n28146_o;
  wire [30:0] n28148_o;
  wire [31:0] n28149_o;
  wire n28151_o;
  wire n28153_o;
  wire n28154_o;
  wire [30:0] n28156_o;
  wire [31:0] n28157_o;
  wire n28159_o;
  wire n28161_o;
  wire n28162_o;
  wire [30:0] n28164_o;
  wire [31:0] n28165_o;
  wire n28167_o;
  wire n28169_o;
  wire n28170_o;
  wire [30:0] n28172_o;
  wire [31:0] n28173_o;
  wire n28175_o;
  wire n28177_o;
  wire n28178_o;
  wire [30:0] n28180_o;
  wire [31:0] n28181_o;
  wire n28183_o;
  wire n28185_o;
  wire n28186_o;
  wire [30:0] n28188_o;
  wire [31:0] n28189_o;
  wire n28191_o;
  wire n28193_o;
  wire n28194_o;
  wire [30:0] n28196_o;
  wire [31:0] n28197_o;
  wire n28199_o;
  wire n28201_o;
  wire n28202_o;
  wire [30:0] n28204_o;
  wire [31:0] n28205_o;
  wire n28207_o;
  wire n28209_o;
  wire n28210_o;
  wire [30:0] n28212_o;
  wire [31:0] n28213_o;
  wire n28215_o;
  wire n28217_o;
  wire n28218_o;
  wire [30:0] n28220_o;
  wire [31:0] n28221_o;
  wire n28223_o;
  wire n28225_o;
  wire n28226_o;
  wire [30:0] n28228_o;
  wire [31:0] n28229_o;
  wire n28231_o;
  wire n28233_o;
  wire n28234_o;
  wire [30:0] n28236_o;
  wire [31:0] n28237_o;
  wire n28239_o;
  wire n28241_o;
  wire n28242_o;
  wire [30:0] n28244_o;
  wire [31:0] n28245_o;
  wire n28247_o;
  wire n28249_o;
  wire n28250_o;
  wire [30:0] n28252_o;
  wire [31:0] n28253_o;
  wire n28255_o;
  wire n28257_o;
  wire n28258_o;
  wire [30:0] n28260_o;
  wire [31:0] n28261_o;
  wire n28263_o;
  wire n28265_o;
  wire n28266_o;
  wire [30:0] n28268_o;
  wire [31:0] n28269_o;
  wire n28271_o;
  wire n28273_o;
  wire n28274_o;
  wire [30:0] n28276_o;
  wire [31:0] n28277_o;
  wire n28279_o;
  wire n28281_o;
  wire n28282_o;
  wire [30:0] n28284_o;
  wire [31:0] n28285_o;
  wire n28287_o;
  wire n28289_o;
  wire n28290_o;
  wire [30:0] n28292_o;
  wire [31:0] n28293_o;
  wire n28295_o;
  wire n28297_o;
  wire n28298_o;
  wire [30:0] n28300_o;
  wire [31:0] n28301_o;
  wire n28303_o;
  wire n28305_o;
  wire n28306_o;
  wire [30:0] n28308_o;
  wire [31:0] n28309_o;
  wire n28311_o;
  wire n28313_o;
  wire n28314_o;
  wire [30:0] n28316_o;
  wire [31:0] n28317_o;
  wire n28319_o;
  wire n28321_o;
  wire n28322_o;
  wire [30:0] n28324_o;
  wire [31:0] n28325_o;
  wire n28327_o;
  wire n28329_o;
  wire n28330_o;
  wire [30:0] n28332_o;
  wire [31:0] n28333_o;
  wire n28335_o;
  wire n28337_o;
  wire n28338_o;
  wire [30:0] n28340_o;
  wire [31:0] n28341_o;
  wire n28343_o;
  wire n28345_o;
  wire n28346_o;
  wire [30:0] n28348_o;
  wire [31:0] n28349_o;
  wire n28351_o;
  wire n28353_o;
  wire n28354_o;
  wire [30:0] n28356_o;
  wire [31:0] n28357_o;
  wire n28359_o;
  wire n28361_o;
  wire n28362_o;
  wire [30:0] n28364_o;
  wire [31:0] n28365_o;
  wire n28367_o;
  wire n28369_o;
  wire n28370_o;
  wire [30:0] n28372_o;
  wire [31:0] n28373_o;
  wire n28375_o;
  wire n28377_o;
  wire n28378_o;
  wire [30:0] n28380_o;
  wire [31:0] n28381_o;
  wire n28383_o;
  wire n28385_o;
  wire n28386_o;
  wire [30:0] n28388_o;
  wire [31:0] n28389_o;
  wire n28391_o;
  wire n28393_o;
  wire n28394_o;
  wire n28395_o;
  wire [30:0] n28396_o;
  wire [31:0] n28397_o;
  wire n28399_o;
  wire n28401_o;
  wire [63:0] n28402_o;
  wire n28409_o;
  wire n28410_o;
  wire [30:0] n28411_o;
  wire [31:0] n28412_o;
  wire n28414_o;
  wire n28417_o;
  wire [30:0] n28418_o;
  wire [31:0] n28419_o;
  wire n28421_o;
  wire n28424_o;
  wire [30:0] n28425_o;
  wire [31:0] n28426_o;
  wire n28428_o;
  wire n28431_o;
  wire [30:0] n28432_o;
  wire [31:0] n28433_o;
  wire n28435_o;
  wire n28438_o;
  wire [30:0] n28439_o;
  wire [31:0] n28440_o;
  wire n28442_o;
  wire n28445_o;
  wire [30:0] n28446_o;
  wire [31:0] n28447_o;
  wire n28449_o;
  wire n28452_o;
  wire [30:0] n28453_o;
  wire [31:0] n28454_o;
  wire n28456_o;
  wire n28459_o;
  wire [30:0] n28460_o;
  wire [31:0] n28461_o;
  wire n28463_o;
  wire n28466_o;
  wire [30:0] n28467_o;
  wire [31:0] n28468_o;
  wire n28470_o;
  wire n28473_o;
  wire [30:0] n28474_o;
  wire [31:0] n28475_o;
  wire n28477_o;
  wire n28480_o;
  wire [30:0] n28481_o;
  wire [31:0] n28482_o;
  wire n28484_o;
  wire n28487_o;
  wire [30:0] n28488_o;
  wire [31:0] n28489_o;
  wire n28491_o;
  wire n28494_o;
  wire [30:0] n28495_o;
  wire [31:0] n28496_o;
  wire n28498_o;
  wire n28501_o;
  wire [30:0] n28502_o;
  wire [31:0] n28503_o;
  wire n28505_o;
  wire n28508_o;
  wire [30:0] n28509_o;
  wire [31:0] n28510_o;
  wire n28512_o;
  wire n28515_o;
  wire [30:0] n28516_o;
  wire [31:0] n28517_o;
  wire n28519_o;
  wire n28522_o;
  wire [30:0] n28523_o;
  wire [31:0] n28524_o;
  wire n28526_o;
  wire n28529_o;
  wire [30:0] n28530_o;
  wire [31:0] n28531_o;
  wire n28533_o;
  wire n28536_o;
  wire [30:0] n28537_o;
  wire [31:0] n28538_o;
  wire n28540_o;
  wire n28543_o;
  wire [30:0] n28544_o;
  wire [31:0] n28545_o;
  wire n28547_o;
  wire n28550_o;
  wire [30:0] n28551_o;
  wire [31:0] n28552_o;
  wire n28554_o;
  wire n28557_o;
  wire [30:0] n28558_o;
  wire [31:0] n28559_o;
  wire n28561_o;
  wire n28564_o;
  wire [30:0] n28565_o;
  wire [31:0] n28566_o;
  wire n28568_o;
  wire n28571_o;
  wire [30:0] n28572_o;
  wire [31:0] n28573_o;
  wire n28575_o;
  wire n28578_o;
  wire [30:0] n28579_o;
  wire [31:0] n28580_o;
  wire n28582_o;
  wire n28585_o;
  wire [30:0] n28586_o;
  wire [31:0] n28587_o;
  wire n28589_o;
  wire n28592_o;
  wire [30:0] n28593_o;
  wire [31:0] n28594_o;
  wire n28596_o;
  wire n28599_o;
  wire [30:0] n28600_o;
  wire [31:0] n28601_o;
  wire n28603_o;
  wire n28606_o;
  wire [30:0] n28607_o;
  wire [31:0] n28608_o;
  wire n28610_o;
  wire n28613_o;
  wire [30:0] n28614_o;
  wire [31:0] n28615_o;
  wire n28617_o;
  wire n28620_o;
  wire [30:0] n28621_o;
  wire [31:0] n28622_o;
  wire n28624_o;
  wire n28627_o;
  wire [30:0] n28628_o;
  wire [31:0] n28629_o;
  wire n28631_o;
  wire n28634_o;
  wire [30:0] n28635_o;
  wire [31:0] n28636_o;
  wire n28638_o;
  wire n28641_o;
  wire [30:0] n28642_o;
  wire [31:0] n28643_o;
  wire n28645_o;
  wire n28648_o;
  wire [30:0] n28649_o;
  wire [31:0] n28650_o;
  wire n28652_o;
  wire n28655_o;
  wire [30:0] n28656_o;
  wire [31:0] n28657_o;
  wire n28659_o;
  wire n28662_o;
  wire [30:0] n28663_o;
  wire [31:0] n28664_o;
  wire n28666_o;
  wire n28669_o;
  wire [30:0] n28670_o;
  wire [31:0] n28671_o;
  wire n28673_o;
  wire n28676_o;
  wire [30:0] n28677_o;
  wire [31:0] n28678_o;
  wire n28680_o;
  wire n28683_o;
  wire [30:0] n28684_o;
  wire [31:0] n28685_o;
  wire n28687_o;
  wire n28690_o;
  wire [30:0] n28691_o;
  wire [31:0] n28692_o;
  wire n28694_o;
  wire n28697_o;
  wire [30:0] n28698_o;
  wire [31:0] n28699_o;
  wire n28701_o;
  wire n28704_o;
  wire [30:0] n28705_o;
  wire [31:0] n28706_o;
  wire n28708_o;
  wire n28711_o;
  wire [30:0] n28712_o;
  wire [31:0] n28713_o;
  wire n28715_o;
  wire n28718_o;
  wire [30:0] n28719_o;
  wire [31:0] n28720_o;
  wire n28722_o;
  wire n28725_o;
  wire [30:0] n28726_o;
  wire [31:0] n28727_o;
  wire n28729_o;
  wire n28732_o;
  wire [30:0] n28733_o;
  wire [31:0] n28734_o;
  wire n28736_o;
  wire n28739_o;
  wire [30:0] n28740_o;
  wire [31:0] n28741_o;
  wire n28743_o;
  wire n28746_o;
  wire [30:0] n28747_o;
  wire [31:0] n28748_o;
  wire n28750_o;
  wire n28753_o;
  wire [30:0] n28754_o;
  wire [31:0] n28755_o;
  wire n28757_o;
  wire n28760_o;
  wire [30:0] n28761_o;
  wire [31:0] n28762_o;
  wire n28764_o;
  wire n28767_o;
  wire [30:0] n28768_o;
  wire [31:0] n28769_o;
  wire n28771_o;
  wire n28774_o;
  wire [30:0] n28775_o;
  wire [31:0] n28776_o;
  wire n28778_o;
  wire n28781_o;
  wire [30:0] n28782_o;
  wire [31:0] n28783_o;
  wire n28785_o;
  wire n28788_o;
  wire [30:0] n28789_o;
  wire [31:0] n28790_o;
  wire n28792_o;
  wire n28795_o;
  wire [30:0] n28796_o;
  wire [31:0] n28797_o;
  wire n28799_o;
  wire n28802_o;
  wire [30:0] n28803_o;
  wire [31:0] n28804_o;
  wire n28806_o;
  wire n28809_o;
  wire [30:0] n28810_o;
  wire [31:0] n28811_o;
  wire n28813_o;
  wire n28816_o;
  wire [30:0] n28817_o;
  wire [31:0] n28818_o;
  wire n28820_o;
  wire n28823_o;
  wire [30:0] n28824_o;
  wire [31:0] n28825_o;
  wire n28827_o;
  wire n28830_o;
  wire [30:0] n28831_o;
  wire [31:0] n28832_o;
  wire n28834_o;
  wire n28837_o;
  wire [30:0] n28838_o;
  wire [31:0] n28839_o;
  wire n28841_o;
  wire n28844_o;
  wire [30:0] n28845_o;
  wire [31:0] n28846_o;
  wire n28848_o;
  wire n28851_o;
  wire [30:0] n28852_o;
  wire [31:0] n28853_o;
  wire n28855_o;
  wire n28858_o;
  wire [63:0] n28859_o;
  wire [63:0] n28861_o;
  wire n28863_o;
  wire n28864_o;
  wire n28865_o;
  wire n28867_o;
  wire n28868_o;
  wire [5:0] n28870_o;
  wire [5:0] n28871_o;
  wire n28872_o;
  wire n28873_o;
  wire n28876_o;
  wire [1:0] n28877_o;
  wire [1:0] n28878_o;
  wire [1:0] n28879_o;
  wire [63:0] n28880_o;
  wire [63:0] n28881_o;
  wire [63:0] n28882_o;
  wire [63:0] n28883_o;
  wire [63:0] n28884_o;
  wire [63:0] n28885_o;
  wire n28887_o;
  wire [63:0] n28888_o;
  wire [63:0] n28889_o;
  wire [63:0] n28890_o;
  wire [63:0] n28891_o;
  wire [63:0] n28892_o;
  wire [63:0] n28893_o;
  wire n28895_o;
  wire [63:0] n28896_o;
  wire n28898_o;
  wire [63:0] n28899_o;
  wire [63:0] n28900_o;
  wire [2:0] n28901_o;
  reg [63:0] n28902_o;
  wire n28904_o;
  wire [63:0] n28905_o;
  wire [63:0] n28906_o;
  wire n28907_o;
  wire n28909_o;
  assign result = n28902_o;
  assign carry_out = n28909_o;
  /* rotator.vhdl:25:12  */
  assign repl32 = n27782_o; // (signal)
  /* rotator.vhdl:26:12  */
  assign rot_count = n27786_o; // (signal)
  /* rotator.vhdl:27:12  */
  assign rot1 = n27804_o; // (signal)
  /* rotator.vhdl:27:18  */
  assign rot2 = n27822_o; // (signal)
  /* rotator.vhdl:27:24  */
  assign rot = n27840_o; // (signal)
  /* rotator.vhdl:28:12  */
  assign sh = n27845_o; // (signal)
  /* rotator.vhdl:28:16  */
  assign mb = n27867_o; // (signal)
  /* rotator.vhdl:28:20  */
  assign me = n27884_o; // (signal)
  /* rotator.vhdl:29:12  */
  assign mr = n28402_o; // (signal)
  /* rotator.vhdl:29:16  */
  assign ml = n28861_o; // (signal)
  /* rotator.vhdl:30:12  */
  assign output_mode = n28879_o; // (signal)
  /* rotator.vhdl:65:23  */
  assign n27734_o = rs[31:0];
  /* rotator.vhdl:68:34  */
  assign n27735_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27736_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27737_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27738_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27739_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27740_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27741_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27742_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27743_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27744_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27745_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27746_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27747_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27748_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27749_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27750_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27751_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27752_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27753_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27754_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27755_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27756_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27757_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27758_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27759_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27760_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27761_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27762_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27763_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27764_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27765_o = rs[31];
  /* rotator.vhdl:68:34  */
  assign n27766_o = rs[31];
  /* common.vhdl:175:14  */
  assign n27767_o = {n27735_o, n27736_o, n27737_o, n27738_o};
  /* common.vhdl:175:14  */
  assign n27768_o = {n27739_o, n27740_o, n27741_o, n27742_o};
  /* common.vhdl:175:14  */
  assign n27769_o = {n27743_o, n27744_o, n27745_o, n27746_o};
  assign n27770_o = {n27747_o, n27748_o, n27749_o, n27750_o};
  /* common.vhdl:175:14  */
  assign n27771_o = {n27751_o, n27752_o, n27753_o, n27754_o};
  assign n27772_o = {n27755_o, n27756_o, n27757_o, n27758_o};
  /* common.vhdl:175:14  */
  assign n27773_o = {n27759_o, n27760_o, n27761_o, n27762_o};
  /* common.vhdl:175:14  */
  assign n27774_o = {n27763_o, n27764_o, n27765_o, n27766_o};
  assign n27775_o = {n27767_o, n27768_o, n27769_o, n27770_o};
  /* common.vhdl:175:14  */
  assign n27776_o = {n27771_o, n27772_o, n27773_o, n27774_o};
  assign n27777_o = {n27775_o, n27776_o};
  /* rotator.vhdl:70:23  */
  assign n27778_o = rs[63:32];
  /* rotator.vhdl:66:9  */
  assign n27779_o = sign_ext_rs ? n27777_o : n27778_o;
  /* rotator.vhdl:64:9  */
  assign n27780_o = is_32bit ? n27734_o : n27779_o;
  /* rotator.vhdl:72:28  */
  assign n27781_o = rs[31:0];
  /* rotator.vhdl:72:24  */
  assign n27782_o = {n27780_o, n27781_o};
  /* rotator.vhdl:76:58  */
  assign n27783_o = shift[5:0];
  /* rotator.vhdl:76:44  */
  assign n27784_o = -n27783_o;
  /* rotator.vhdl:78:31  */
  assign n27785_o = shift[5:0];
  /* rotator.vhdl:75:9  */
  assign n27786_o = right_shift ? n27784_o : n27785_o;
  /* rotator.vhdl:87:23  */
  assign n27787_o = rot_count[1:0];
  /* rotator.vhdl:88:13  */
  assign n27789_o = n27787_o == 2'b00;
  /* rotator.vhdl:91:31  */
  assign n27790_o = repl32[62:0];
  /* rotator.vhdl:91:53  */
  assign n27791_o = repl32[63];
  /* rotator.vhdl:91:45  */
  assign n27792_o = {n27790_o, n27791_o};
  /* rotator.vhdl:90:13  */
  assign n27794_o = n27787_o == 2'b01;
  /* rotator.vhdl:93:31  */
  assign n27795_o = repl32[61:0];
  /* rotator.vhdl:93:53  */
  assign n27796_o = repl32[63:62];
  /* rotator.vhdl:93:45  */
  assign n27797_o = {n27795_o, n27796_o};
  /* rotator.vhdl:92:13  */
  assign n27799_o = n27787_o == 2'b10;
  /* rotator.vhdl:95:31  */
  assign n27800_o = repl32[60:0];
  /* rotator.vhdl:95:53  */
  assign n27801_o = repl32[63:61];
  /* rotator.vhdl:95:45  */
  assign n27802_o = {n27800_o, n27801_o};
  assign n27803_o = {n27799_o, n27794_o, n27789_o};
  /* rotator.vhdl:87:9  */
  always @*
    case (n27803_o)
      3'b100: n27804_o = n27797_o;
      3'b010: n27804_o = n27792_o;
      3'b001: n27804_o = repl32;
      default: n27804_o = n27802_o;
    endcase
  /* rotator.vhdl:98:23  */
  assign n27805_o = rot_count[3:2];
  /* rotator.vhdl:99:13  */
  assign n27807_o = n27805_o == 2'b00;
  /* rotator.vhdl:102:29  */
  assign n27808_o = rot1[59:0];
  /* rotator.vhdl:102:49  */
  assign n27809_o = rot1[63:60];
  /* rotator.vhdl:102:43  */
  assign n27810_o = {n27808_o, n27809_o};
  /* rotator.vhdl:101:13  */
  assign n27812_o = n27805_o == 2'b01;
  /* rotator.vhdl:104:29  */
  assign n27813_o = rot1[55:0];
  /* rotator.vhdl:104:49  */
  assign n27814_o = rot1[63:56];
  /* rotator.vhdl:104:43  */
  assign n27815_o = {n27813_o, n27814_o};
  /* rotator.vhdl:103:13  */
  assign n27817_o = n27805_o == 2'b10;
  /* rotator.vhdl:106:29  */
  assign n27818_o = rot1[51:0];
  /* rotator.vhdl:106:49  */
  assign n27819_o = rot1[63:52];
  /* rotator.vhdl:106:43  */
  assign n27820_o = {n27818_o, n27819_o};
  /* control.vhdl:109:65  */
  assign n27821_o = {n27817_o, n27812_o, n27807_o};
  /* rotator.vhdl:98:9  */
  always @*
    case (n27821_o)
      3'b100: n27822_o = n27815_o;
      3'b010: n27822_o = n27810_o;
      3'b001: n27822_o = rot1;
      default: n27822_o = n27820_o;
    endcase
  /* rotator.vhdl:109:23  */
  assign n27823_o = rot_count[5:4];
  /* rotator.vhdl:110:13  */
  assign n27825_o = n27823_o == 2'b00;
  /* rotator.vhdl:113:28  */
  assign n27826_o = rot2[47:0];
  /* rotator.vhdl:113:48  */
  assign n27827_o = rot2[63:48];
  /* rotator.vhdl:113:42  */
  assign n27828_o = {n27826_o, n27827_o};
  /* rotator.vhdl:112:13  */
  assign n27830_o = n27823_o == 2'b01;
  /* rotator.vhdl:115:28  */
  assign n27831_o = rot2[31:0];
  /* rotator.vhdl:115:48  */
  assign n27832_o = rot2[63:32];
  /* rotator.vhdl:115:42  */
  assign n27833_o = {n27831_o, n27832_o};
  /* rotator.vhdl:114:13  */
  assign n27835_o = n27823_o == 2'b10;
  /* rotator.vhdl:117:28  */
  assign n27836_o = rot2[15:0];
  /* rotator.vhdl:117:48  */
  assign n27837_o = rot2[63:16];
  /* rotator.vhdl:117:42  */
  assign n27838_o = {n27836_o, n27837_o};
  assign n27839_o = {n27835_o, n27830_o, n27825_o};
  /* rotator.vhdl:109:9  */
  always @*
    case (n27839_o)
      3'b100: n27840_o = n27833_o;
      3'b010: n27840_o = n27828_o;
      3'b001: n27840_o = rot2;
      default: n27840_o = n27838_o;
    endcase
  /* rotator.vhdl:121:21  */
  assign n27841_o = shift[6];
  /* rotator.vhdl:121:29  */
  assign n27842_o = ~is_32bit;
  /* rotator.vhdl:121:25  */
  assign n27843_o = n27841_o & n27842_o;
  /* rotator.vhdl:121:50  */
  assign n27844_o = shift[5:0];
  /* rotator.vhdl:121:43  */
  assign n27845_o = {n27843_o, n27844_o};
  /* rotator.vhdl:126:34  */
  assign n27846_o = insn[10:6];
  /* rotator.vhdl:126:28  */
  assign n27848_o = {2'b01, n27846_o};
  /* rotator.vhdl:128:33  */
  assign n27849_o = insn[5];
  /* rotator.vhdl:128:27  */
  assign n27851_o = {1'b0, n27849_o};
  /* rotator.vhdl:128:43  */
  assign n27852_o = insn[10:6];
  /* rotator.vhdl:128:37  */
  assign n27853_o = {n27851_o, n27852_o};
  /* rotator.vhdl:125:13  */
  assign n27854_o = is_32bit ? n27848_o : n27853_o;
  /* rotator.vhdl:133:25  */
  assign n27855_o = sh[5];
  /* rotator.vhdl:133:37  */
  assign n27856_o = sh[5];
  /* rotator.vhdl:133:31  */
  assign n27857_o = ~n27856_o;
  /* rotator.vhdl:133:29  */
  assign n27858_o = {n27855_o, n27857_o};
  /* rotator.vhdl:133:45  */
  assign n27859_o = sh[4:0];
  /* rotator.vhdl:133:41  */
  assign n27860_o = {n27858_o, n27859_o};
  /* rotator.vhdl:132:13  */
  assign n27861_o = is_32bit ? n27860_o : sh;
  /* rotator.vhdl:138:24  */
  assign n27863_o = {1'b0, is_32bit};
  /* rotator.vhdl:138:35  */
  assign n27865_o = {n27863_o, 5'b00000};
  /* rotator.vhdl:130:9  */
  assign n27866_o = right_shift ? n27861_o : n27865_o;
  /* rotator.vhdl:124:9  */
  assign n27867_o = clear_left ? n27854_o : n27866_o;
  /* rotator.vhdl:140:30  */
  assign n27868_o = clear_right & is_32bit;
  /* rotator.vhdl:141:30  */
  assign n27869_o = insn[5:1];
  /* rotator.vhdl:141:24  */
  assign n27871_o = {2'b01, n27869_o};
  /* rotator.vhdl:142:48  */
  assign n27872_o = ~clear_left;
  /* rotator.vhdl:142:33  */
  assign n27873_o = clear_right & n27872_o;
  /* rotator.vhdl:143:29  */
  assign n27874_o = insn[5];
  /* rotator.vhdl:143:23  */
  assign n27876_o = {1'b0, n27874_o};
  /* rotator.vhdl:143:39  */
  assign n27877_o = insn[10:6];
  /* rotator.vhdl:143:33  */
  assign n27878_o = {n27876_o, n27877_o};
  /* rotator.vhdl:146:21  */
  assign n27879_o = sh[6];
  /* rotator.vhdl:146:33  */
  assign n27880_o = sh[5:0];
  /* rotator.vhdl:146:27  */
  assign n27881_o = ~n27880_o;
  /* rotator.vhdl:146:25  */
  assign n27882_o = {n27879_o, n27881_o};
  /* rotator.vhdl:142:9  */
  assign n27883_o = n27873_o ? n27878_o : n27882_o;
  /* rotator.vhdl:140:9  */
  assign n27884_o = n27868_o ? n27871_o : n27883_o;
  /* rotator.vhdl:38:21  */
  assign n27891_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27892_o = {1'b0, n27891_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27894_o = $signed(32'b00000000000000000000000000000000) >= $signed(n27892_o);
  /* rotator.vhdl:38:13  */
  assign n27897_o = n27894_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:38:21  */
  assign n27900_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27901_o = {1'b0, n27900_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27903_o = $signed(32'b00000000000000000000000000000001) >= $signed(n27901_o);
  assign n27905_o = n27898_o[62];
  /* rotator.vhdl:38:13  */
  assign n27906_o = n27903_o ? 1'b1 : n27905_o;
  /* rotator.vhdl:38:21  */
  assign n27908_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27909_o = {1'b0, n27908_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27911_o = $signed(32'b00000000000000000000000000000010) >= $signed(n27909_o);
  assign n27913_o = n27898_o[61];
  /* rotator.vhdl:38:13  */
  assign n27914_o = n27911_o ? 1'b1 : n27913_o;
  /* rotator.vhdl:38:21  */
  assign n27916_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27917_o = {1'b0, n27916_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27919_o = $signed(32'b00000000000000000000000000000011) >= $signed(n27917_o);
  assign n27921_o = n27898_o[60];
  /* rotator.vhdl:38:13  */
  assign n27922_o = n27919_o ? 1'b1 : n27921_o;
  /* rotator.vhdl:38:21  */
  assign n27924_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27925_o = {1'b0, n27924_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27927_o = $signed(32'b00000000000000000000000000000100) >= $signed(n27925_o);
  assign n27929_o = n27898_o[59];
  /* rotator.vhdl:38:13  */
  assign n27930_o = n27927_o ? 1'b1 : n27929_o;
  /* rotator.vhdl:38:21  */
  assign n27932_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27933_o = {1'b0, n27932_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27935_o = $signed(32'b00000000000000000000000000000101) >= $signed(n27933_o);
  assign n27937_o = n27898_o[58];
  /* rotator.vhdl:38:13  */
  assign n27938_o = n27935_o ? 1'b1 : n27937_o;
  /* rotator.vhdl:38:21  */
  assign n27940_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27941_o = {1'b0, n27940_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27943_o = $signed(32'b00000000000000000000000000000110) >= $signed(n27941_o);
  assign n27945_o = n27898_o[57];
  /* rotator.vhdl:38:13  */
  assign n27946_o = n27943_o ? 1'b1 : n27945_o;
  /* rotator.vhdl:38:21  */
  assign n27948_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27949_o = {1'b0, n27948_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27951_o = $signed(32'b00000000000000000000000000000111) >= $signed(n27949_o);
  assign n27953_o = n27898_o[56];
  /* rotator.vhdl:38:13  */
  assign n27954_o = n27951_o ? 1'b1 : n27953_o;
  /* rotator.vhdl:38:21  */
  assign n27956_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27957_o = {1'b0, n27956_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27959_o = $signed(32'b00000000000000000000000000001000) >= $signed(n27957_o);
  assign n27961_o = n27898_o[55];
  /* rotator.vhdl:38:13  */
  assign n27962_o = n27959_o ? 1'b1 : n27961_o;
  /* rotator.vhdl:38:21  */
  assign n27964_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27965_o = {1'b0, n27964_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27967_o = $signed(32'b00000000000000000000000000001001) >= $signed(n27965_o);
  assign n27969_o = n27898_o[54];
  /* rotator.vhdl:38:13  */
  assign n27970_o = n27967_o ? 1'b1 : n27969_o;
  /* rotator.vhdl:38:21  */
  assign n27972_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27973_o = {1'b0, n27972_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27975_o = $signed(32'b00000000000000000000000000001010) >= $signed(n27973_o);
  assign n27977_o = n27898_o[53];
  /* rotator.vhdl:38:13  */
  assign n27978_o = n27975_o ? 1'b1 : n27977_o;
  /* rotator.vhdl:38:21  */
  assign n27980_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27981_o = {1'b0, n27980_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27983_o = $signed(32'b00000000000000000000000000001011) >= $signed(n27981_o);
  assign n27985_o = n27898_o[52];
  /* rotator.vhdl:38:13  */
  assign n27986_o = n27983_o ? 1'b1 : n27985_o;
  /* rotator.vhdl:38:21  */
  assign n27988_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27989_o = {1'b0, n27988_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27991_o = $signed(32'b00000000000000000000000000001100) >= $signed(n27989_o);
  assign n27993_o = n27898_o[51];
  /* rotator.vhdl:38:13  */
  assign n27994_o = n27991_o ? 1'b1 : n27993_o;
  /* rotator.vhdl:38:21  */
  assign n27996_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27997_o = {1'b0, n27996_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n27999_o = $signed(32'b00000000000000000000000000001101) >= $signed(n27997_o);
  assign n28001_o = n27898_o[50];
  /* rotator.vhdl:38:13  */
  assign n28002_o = n27999_o ? 1'b1 : n28001_o;
  /* rotator.vhdl:38:21  */
  assign n28004_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28005_o = {1'b0, n28004_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28007_o = $signed(32'b00000000000000000000000000001110) >= $signed(n28005_o);
  assign n28009_o = n27898_o[49];
  /* rotator.vhdl:38:13  */
  assign n28010_o = n28007_o ? 1'b1 : n28009_o;
  /* rotator.vhdl:38:21  */
  assign n28012_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28013_o = {1'b0, n28012_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28015_o = $signed(32'b00000000000000000000000000001111) >= $signed(n28013_o);
  assign n28017_o = n27898_o[48];
  /* rotator.vhdl:38:13  */
  assign n28018_o = n28015_o ? 1'b1 : n28017_o;
  /* rotator.vhdl:38:21  */
  assign n28020_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28021_o = {1'b0, n28020_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28023_o = $signed(32'b00000000000000000000000000010000) >= $signed(n28021_o);
  assign n28025_o = n27898_o[47];
  /* rotator.vhdl:38:13  */
  assign n28026_o = n28023_o ? 1'b1 : n28025_o;
  /* rotator.vhdl:38:21  */
  assign n28028_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28029_o = {1'b0, n28028_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28031_o = $signed(32'b00000000000000000000000000010001) >= $signed(n28029_o);
  assign n28033_o = n27898_o[46];
  /* rotator.vhdl:38:13  */
  assign n28034_o = n28031_o ? 1'b1 : n28033_o;
  /* rotator.vhdl:38:21  */
  assign n28036_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28037_o = {1'b0, n28036_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28039_o = $signed(32'b00000000000000000000000000010010) >= $signed(n28037_o);
  assign n28041_o = n27898_o[45];
  /* rotator.vhdl:38:13  */
  assign n28042_o = n28039_o ? 1'b1 : n28041_o;
  /* rotator.vhdl:38:21  */
  assign n28044_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28045_o = {1'b0, n28044_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28047_o = $signed(32'b00000000000000000000000000010011) >= $signed(n28045_o);
  assign n28049_o = n27898_o[44];
  /* rotator.vhdl:38:13  */
  assign n28050_o = n28047_o ? 1'b1 : n28049_o;
  /* rotator.vhdl:38:21  */
  assign n28052_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28053_o = {1'b0, n28052_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28055_o = $signed(32'b00000000000000000000000000010100) >= $signed(n28053_o);
  assign n28057_o = n27898_o[43];
  /* rotator.vhdl:38:13  */
  assign n28058_o = n28055_o ? 1'b1 : n28057_o;
  /* rotator.vhdl:38:21  */
  assign n28060_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28061_o = {1'b0, n28060_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28063_o = $signed(32'b00000000000000000000000000010101) >= $signed(n28061_o);
  assign n28065_o = n27898_o[42];
  /* rotator.vhdl:38:13  */
  assign n28066_o = n28063_o ? 1'b1 : n28065_o;
  /* rotator.vhdl:38:21  */
  assign n28068_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28069_o = {1'b0, n28068_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28071_o = $signed(32'b00000000000000000000000000010110) >= $signed(n28069_o);
  assign n28073_o = n27898_o[41];
  /* rotator.vhdl:38:13  */
  assign n28074_o = n28071_o ? 1'b1 : n28073_o;
  /* rotator.vhdl:38:21  */
  assign n28076_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28077_o = {1'b0, n28076_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28079_o = $signed(32'b00000000000000000000000000010111) >= $signed(n28077_o);
  assign n28081_o = n27898_o[40];
  /* rotator.vhdl:38:13  */
  assign n28082_o = n28079_o ? 1'b1 : n28081_o;
  /* rotator.vhdl:38:21  */
  assign n28084_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28085_o = {1'b0, n28084_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28087_o = $signed(32'b00000000000000000000000000011000) >= $signed(n28085_o);
  assign n28089_o = n27898_o[39];
  /* rotator.vhdl:38:13  */
  assign n28090_o = n28087_o ? 1'b1 : n28089_o;
  /* rotator.vhdl:38:21  */
  assign n28092_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28093_o = {1'b0, n28092_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28095_o = $signed(32'b00000000000000000000000000011001) >= $signed(n28093_o);
  assign n28097_o = n27898_o[38];
  /* rotator.vhdl:38:13  */
  assign n28098_o = n28095_o ? 1'b1 : n28097_o;
  /* rotator.vhdl:38:21  */
  assign n28100_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28101_o = {1'b0, n28100_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28103_o = $signed(32'b00000000000000000000000000011010) >= $signed(n28101_o);
  assign n28105_o = n27898_o[37];
  /* rotator.vhdl:38:13  */
  assign n28106_o = n28103_o ? 1'b1 : n28105_o;
  /* rotator.vhdl:38:21  */
  assign n28108_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28109_o = {1'b0, n28108_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28111_o = $signed(32'b00000000000000000000000000011011) >= $signed(n28109_o);
  assign n28113_o = n27898_o[36];
  /* rotator.vhdl:38:13  */
  assign n28114_o = n28111_o ? 1'b1 : n28113_o;
  /* rotator.vhdl:38:21  */
  assign n28116_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28117_o = {1'b0, n28116_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28119_o = $signed(32'b00000000000000000000000000011100) >= $signed(n28117_o);
  assign n28121_o = n27898_o[35];
  /* rotator.vhdl:38:13  */
  assign n28122_o = n28119_o ? 1'b1 : n28121_o;
  /* rotator.vhdl:38:21  */
  assign n28124_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28125_o = {1'b0, n28124_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28127_o = $signed(32'b00000000000000000000000000011101) >= $signed(n28125_o);
  assign n28129_o = n27898_o[34];
  /* rotator.vhdl:38:13  */
  assign n28130_o = n28127_o ? 1'b1 : n28129_o;
  /* rotator.vhdl:38:21  */
  assign n28132_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28133_o = {1'b0, n28132_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28135_o = $signed(32'b00000000000000000000000000011110) >= $signed(n28133_o);
  assign n28137_o = n27898_o[33];
  /* rotator.vhdl:38:13  */
  assign n28138_o = n28135_o ? 1'b1 : n28137_o;
  /* rotator.vhdl:38:21  */
  assign n28140_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28141_o = {1'b0, n28140_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28143_o = $signed(32'b00000000000000000000000000011111) >= $signed(n28141_o);
  assign n28145_o = n27898_o[32];
  /* rotator.vhdl:38:13  */
  assign n28146_o = n28143_o ? 1'b1 : n28145_o;
  /* rotator.vhdl:38:21  */
  assign n28148_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28149_o = {1'b0, n28148_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28151_o = $signed(32'b00000000000000000000000000100000) >= $signed(n28149_o);
  assign n28153_o = n27898_o[31];
  /* rotator.vhdl:38:13  */
  assign n28154_o = n28151_o ? 1'b1 : n28153_o;
  /* rotator.vhdl:38:21  */
  assign n28156_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28157_o = {1'b0, n28156_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28159_o = $signed(32'b00000000000000000000000000100001) >= $signed(n28157_o);
  assign n28161_o = n27898_o[30];
  /* rotator.vhdl:38:13  */
  assign n28162_o = n28159_o ? 1'b1 : n28161_o;
  /* rotator.vhdl:38:21  */
  assign n28164_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28165_o = {1'b0, n28164_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28167_o = $signed(32'b00000000000000000000000000100010) >= $signed(n28165_o);
  assign n28169_o = n27898_o[29];
  /* rotator.vhdl:38:13  */
  assign n28170_o = n28167_o ? 1'b1 : n28169_o;
  /* rotator.vhdl:38:21  */
  assign n28172_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28173_o = {1'b0, n28172_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28175_o = $signed(32'b00000000000000000000000000100011) >= $signed(n28173_o);
  assign n28177_o = n27898_o[28];
  /* rotator.vhdl:38:13  */
  assign n28178_o = n28175_o ? 1'b1 : n28177_o;
  /* rotator.vhdl:38:21  */
  assign n28180_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28181_o = {1'b0, n28180_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28183_o = $signed(32'b00000000000000000000000000100100) >= $signed(n28181_o);
  assign n28185_o = n27898_o[27];
  /* rotator.vhdl:38:13  */
  assign n28186_o = n28183_o ? 1'b1 : n28185_o;
  /* rotator.vhdl:38:21  */
  assign n28188_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28189_o = {1'b0, n28188_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28191_o = $signed(32'b00000000000000000000000000100101) >= $signed(n28189_o);
  assign n28193_o = n27898_o[26];
  /* rotator.vhdl:38:13  */
  assign n28194_o = n28191_o ? 1'b1 : n28193_o;
  /* rotator.vhdl:38:21  */
  assign n28196_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28197_o = {1'b0, n28196_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28199_o = $signed(32'b00000000000000000000000000100110) >= $signed(n28197_o);
  assign n28201_o = n27898_o[25];
  /* rotator.vhdl:38:13  */
  assign n28202_o = n28199_o ? 1'b1 : n28201_o;
  /* rotator.vhdl:38:21  */
  assign n28204_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28205_o = {1'b0, n28204_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28207_o = $signed(32'b00000000000000000000000000100111) >= $signed(n28205_o);
  assign n28209_o = n27898_o[24];
  /* rotator.vhdl:38:13  */
  assign n28210_o = n28207_o ? 1'b1 : n28209_o;
  /* rotator.vhdl:38:21  */
  assign n28212_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28213_o = {1'b0, n28212_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28215_o = $signed(32'b00000000000000000000000000101000) >= $signed(n28213_o);
  assign n28217_o = n27898_o[23];
  /* rotator.vhdl:38:13  */
  assign n28218_o = n28215_o ? 1'b1 : n28217_o;
  /* rotator.vhdl:38:21  */
  assign n28220_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28221_o = {1'b0, n28220_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28223_o = $signed(32'b00000000000000000000000000101001) >= $signed(n28221_o);
  assign n28225_o = n27898_o[22];
  /* rotator.vhdl:38:13  */
  assign n28226_o = n28223_o ? 1'b1 : n28225_o;
  /* rotator.vhdl:38:21  */
  assign n28228_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28229_o = {1'b0, n28228_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28231_o = $signed(32'b00000000000000000000000000101010) >= $signed(n28229_o);
  assign n28233_o = n27898_o[21];
  /* rotator.vhdl:38:13  */
  assign n28234_o = n28231_o ? 1'b1 : n28233_o;
  /* rotator.vhdl:38:21  */
  assign n28236_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28237_o = {1'b0, n28236_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28239_o = $signed(32'b00000000000000000000000000101011) >= $signed(n28237_o);
  assign n28241_o = n27898_o[20];
  /* rotator.vhdl:38:13  */
  assign n28242_o = n28239_o ? 1'b1 : n28241_o;
  /* rotator.vhdl:38:21  */
  assign n28244_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28245_o = {1'b0, n28244_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28247_o = $signed(32'b00000000000000000000000000101100) >= $signed(n28245_o);
  assign n28249_o = n27898_o[19];
  /* rotator.vhdl:38:13  */
  assign n28250_o = n28247_o ? 1'b1 : n28249_o;
  /* rotator.vhdl:38:21  */
  assign n28252_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28253_o = {1'b0, n28252_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28255_o = $signed(32'b00000000000000000000000000101101) >= $signed(n28253_o);
  assign n28257_o = n27898_o[18];
  /* rotator.vhdl:38:13  */
  assign n28258_o = n28255_o ? 1'b1 : n28257_o;
  /* rotator.vhdl:38:21  */
  assign n28260_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28261_o = {1'b0, n28260_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28263_o = $signed(32'b00000000000000000000000000101110) >= $signed(n28261_o);
  assign n28265_o = n27898_o[17];
  /* rotator.vhdl:38:13  */
  assign n28266_o = n28263_o ? 1'b1 : n28265_o;
  /* rotator.vhdl:38:21  */
  assign n28268_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28269_o = {1'b0, n28268_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28271_o = $signed(32'b00000000000000000000000000101111) >= $signed(n28269_o);
  assign n28273_o = n27898_o[16];
  /* rotator.vhdl:38:13  */
  assign n28274_o = n28271_o ? 1'b1 : n28273_o;
  /* rotator.vhdl:38:21  */
  assign n28276_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28277_o = {1'b0, n28276_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28279_o = $signed(32'b00000000000000000000000000110000) >= $signed(n28277_o);
  assign n28281_o = n27898_o[15];
  /* rotator.vhdl:38:13  */
  assign n28282_o = n28279_o ? 1'b1 : n28281_o;
  /* rotator.vhdl:38:21  */
  assign n28284_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28285_o = {1'b0, n28284_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28287_o = $signed(32'b00000000000000000000000000110001) >= $signed(n28285_o);
  assign n28289_o = n27898_o[14];
  /* rotator.vhdl:38:13  */
  assign n28290_o = n28287_o ? 1'b1 : n28289_o;
  /* rotator.vhdl:38:21  */
  assign n28292_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28293_o = {1'b0, n28292_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28295_o = $signed(32'b00000000000000000000000000110010) >= $signed(n28293_o);
  assign n28297_o = n27898_o[13];
  /* rotator.vhdl:38:13  */
  assign n28298_o = n28295_o ? 1'b1 : n28297_o;
  /* rotator.vhdl:38:21  */
  assign n28300_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28301_o = {1'b0, n28300_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28303_o = $signed(32'b00000000000000000000000000110011) >= $signed(n28301_o);
  assign n28305_o = n27898_o[12];
  /* rotator.vhdl:38:13  */
  assign n28306_o = n28303_o ? 1'b1 : n28305_o;
  /* rotator.vhdl:38:21  */
  assign n28308_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28309_o = {1'b0, n28308_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28311_o = $signed(32'b00000000000000000000000000110100) >= $signed(n28309_o);
  assign n28313_o = n27898_o[11];
  /* rotator.vhdl:38:13  */
  assign n28314_o = n28311_o ? 1'b1 : n28313_o;
  /* rotator.vhdl:38:21  */
  assign n28316_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28317_o = {1'b0, n28316_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28319_o = $signed(32'b00000000000000000000000000110101) >= $signed(n28317_o);
  assign n28321_o = n27898_o[10];
  /* rotator.vhdl:38:13  */
  assign n28322_o = n28319_o ? 1'b1 : n28321_o;
  /* rotator.vhdl:38:21  */
  assign n28324_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28325_o = {1'b0, n28324_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28327_o = $signed(32'b00000000000000000000000000110110) >= $signed(n28325_o);
  assign n28329_o = n27898_o[9];
  /* rotator.vhdl:38:13  */
  assign n28330_o = n28327_o ? 1'b1 : n28329_o;
  /* rotator.vhdl:38:21  */
  assign n28332_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28333_o = {1'b0, n28332_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28335_o = $signed(32'b00000000000000000000000000110111) >= $signed(n28333_o);
  assign n28337_o = n27898_o[8];
  /* rotator.vhdl:38:13  */
  assign n28338_o = n28335_o ? 1'b1 : n28337_o;
  /* rotator.vhdl:38:21  */
  assign n28340_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28341_o = {1'b0, n28340_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28343_o = $signed(32'b00000000000000000000000000111000) >= $signed(n28341_o);
  assign n28345_o = n27898_o[7];
  /* rotator.vhdl:38:13  */
  assign n28346_o = n28343_o ? 1'b1 : n28345_o;
  /* rotator.vhdl:38:21  */
  assign n28348_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28349_o = {1'b0, n28348_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28351_o = $signed(32'b00000000000000000000000000111001) >= $signed(n28349_o);
  assign n28353_o = n27898_o[6];
  /* rotator.vhdl:38:13  */
  assign n28354_o = n28351_o ? 1'b1 : n28353_o;
  /* rotator.vhdl:38:21  */
  assign n28356_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28357_o = {1'b0, n28356_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28359_o = $signed(32'b00000000000000000000000000111010) >= $signed(n28357_o);
  assign n28361_o = n27898_o[5];
  /* rotator.vhdl:38:13  */
  assign n28362_o = n28359_o ? 1'b1 : n28361_o;
  /* rotator.vhdl:38:21  */
  assign n28364_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28365_o = {1'b0, n28364_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28367_o = $signed(32'b00000000000000000000000000111011) >= $signed(n28365_o);
  assign n28369_o = n27898_o[4];
  /* rotator.vhdl:38:13  */
  assign n28370_o = n28367_o ? 1'b1 : n28369_o;
  /* rotator.vhdl:38:21  */
  assign n28372_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28373_o = {1'b0, n28372_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28375_o = $signed(32'b00000000000000000000000000111100) >= $signed(n28373_o);
  assign n28377_o = n27898_o[3];
  /* rotator.vhdl:38:13  */
  assign n28378_o = n28375_o ? 1'b1 : n28377_o;
  /* rotator.vhdl:38:21  */
  assign n28380_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28381_o = {1'b0, n28380_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28383_o = $signed(32'b00000000000000000000000000111101) >= $signed(n28381_o);
  assign n28385_o = n27898_o[2];
  /* rotator.vhdl:38:13  */
  assign n28386_o = n28383_o ? 1'b1 : n28385_o;
  /* rotator.vhdl:38:21  */
  assign n28388_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28389_o = {1'b0, n28388_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28391_o = $signed(32'b00000000000000000000000000111110) >= $signed(n28389_o);
  assign n28393_o = n27898_o[1];
  /* rotator.vhdl:38:13  */
  assign n28394_o = n28391_o ? 1'b1 : n28393_o;
  assign n28395_o = n27898_o[0];
  /* rotator.vhdl:38:21  */
  assign n28396_o = {24'b0, mb};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28397_o = {1'b0, n28396_o};  //  uext
  /* rotator.vhdl:38:18  */
  assign n28399_o = $signed(32'b00000000000000000000000000111111) >= $signed(n28397_o);
  /* rotator.vhdl:38:13  */
  assign n28401_o = n28399_o ? 1'b1 : n28395_o;
  assign n28402_o = {n27897_o, n27906_o, n27914_o, n27922_o, n27930_o, n27938_o, n27946_o, n27954_o, n27962_o, n27970_o, n27978_o, n27986_o, n27994_o, n28002_o, n28010_o, n28018_o, n28026_o, n28034_o, n28042_o, n28050_o, n28058_o, n28066_o, n28074_o, n28082_o, n28090_o, n28098_o, n28106_o, n28114_o, n28122_o, n28130_o, n28138_o, n28146_o, n28154_o, n28162_o, n28170_o, n28178_o, n28186_o, n28194_o, n28202_o, n28210_o, n28218_o, n28226_o, n28234_o, n28242_o, n28250_o, n28258_o, n28266_o, n28274_o, n28282_o, n28290_o, n28298_o, n28306_o, n28314_o, n28322_o, n28330_o, n28338_o, n28346_o, n28354_o, n28362_o, n28370_o, n28378_o, n28386_o, n28394_o, n28401_o};
  /* rotator.vhdl:49:20  */
  assign n28409_o = me[6];
  /* rotator.vhdl:49:24  */
  assign n28410_o = ~n28409_o;
  /* rotator.vhdl:51:25  */
  assign n28411_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28412_o = {1'b0, n28411_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28414_o = $signed(32'b00000000000000000000000000000000) <= $signed(n28412_o);
  /* rotator.vhdl:51:17  */
  assign n28417_o = n28414_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28418_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28419_o = {1'b0, n28418_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28421_o = $signed(32'b00000000000000000000000000000001) <= $signed(n28419_o);
  /* rotator.vhdl:51:17  */
  assign n28424_o = n28421_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28425_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28426_o = {1'b0, n28425_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28428_o = $signed(32'b00000000000000000000000000000010) <= $signed(n28426_o);
  /* rotator.vhdl:51:17  */
  assign n28431_o = n28428_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28432_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28433_o = {1'b0, n28432_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28435_o = $signed(32'b00000000000000000000000000000011) <= $signed(n28433_o);
  /* rotator.vhdl:51:17  */
  assign n28438_o = n28435_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28439_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28440_o = {1'b0, n28439_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28442_o = $signed(32'b00000000000000000000000000000100) <= $signed(n28440_o);
  /* rotator.vhdl:51:17  */
  assign n28445_o = n28442_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28446_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28447_o = {1'b0, n28446_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28449_o = $signed(32'b00000000000000000000000000000101) <= $signed(n28447_o);
  /* rotator.vhdl:51:17  */
  assign n28452_o = n28449_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28453_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28454_o = {1'b0, n28453_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28456_o = $signed(32'b00000000000000000000000000000110) <= $signed(n28454_o);
  /* rotator.vhdl:51:17  */
  assign n28459_o = n28456_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28460_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28461_o = {1'b0, n28460_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28463_o = $signed(32'b00000000000000000000000000000111) <= $signed(n28461_o);
  /* rotator.vhdl:51:17  */
  assign n28466_o = n28463_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28467_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28468_o = {1'b0, n28467_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28470_o = $signed(32'b00000000000000000000000000001000) <= $signed(n28468_o);
  /* rotator.vhdl:51:17  */
  assign n28473_o = n28470_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28474_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28475_o = {1'b0, n28474_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28477_o = $signed(32'b00000000000000000000000000001001) <= $signed(n28475_o);
  /* rotator.vhdl:51:17  */
  assign n28480_o = n28477_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28481_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28482_o = {1'b0, n28481_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28484_o = $signed(32'b00000000000000000000000000001010) <= $signed(n28482_o);
  /* rotator.vhdl:51:17  */
  assign n28487_o = n28484_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28488_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28489_o = {1'b0, n28488_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28491_o = $signed(32'b00000000000000000000000000001011) <= $signed(n28489_o);
  /* rotator.vhdl:51:17  */
  assign n28494_o = n28491_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28495_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28496_o = {1'b0, n28495_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28498_o = $signed(32'b00000000000000000000000000001100) <= $signed(n28496_o);
  /* rotator.vhdl:51:17  */
  assign n28501_o = n28498_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28502_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28503_o = {1'b0, n28502_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28505_o = $signed(32'b00000000000000000000000000001101) <= $signed(n28503_o);
  /* rotator.vhdl:51:17  */
  assign n28508_o = n28505_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28509_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28510_o = {1'b0, n28509_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28512_o = $signed(32'b00000000000000000000000000001110) <= $signed(n28510_o);
  /* rotator.vhdl:51:17  */
  assign n28515_o = n28512_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28516_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28517_o = {1'b0, n28516_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28519_o = $signed(32'b00000000000000000000000000001111) <= $signed(n28517_o);
  /* rotator.vhdl:51:17  */
  assign n28522_o = n28519_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28523_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28524_o = {1'b0, n28523_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28526_o = $signed(32'b00000000000000000000000000010000) <= $signed(n28524_o);
  /* rotator.vhdl:51:17  */
  assign n28529_o = n28526_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28530_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28531_o = {1'b0, n28530_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28533_o = $signed(32'b00000000000000000000000000010001) <= $signed(n28531_o);
  /* rotator.vhdl:51:17  */
  assign n28536_o = n28533_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28537_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28538_o = {1'b0, n28537_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28540_o = $signed(32'b00000000000000000000000000010010) <= $signed(n28538_o);
  /* rotator.vhdl:51:17  */
  assign n28543_o = n28540_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28544_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28545_o = {1'b0, n28544_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28547_o = $signed(32'b00000000000000000000000000010011) <= $signed(n28545_o);
  /* rotator.vhdl:51:17  */
  assign n28550_o = n28547_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28551_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28552_o = {1'b0, n28551_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28554_o = $signed(32'b00000000000000000000000000010100) <= $signed(n28552_o);
  /* rotator.vhdl:51:17  */
  assign n28557_o = n28554_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28558_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28559_o = {1'b0, n28558_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28561_o = $signed(32'b00000000000000000000000000010101) <= $signed(n28559_o);
  /* rotator.vhdl:51:17  */
  assign n28564_o = n28561_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28565_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28566_o = {1'b0, n28565_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28568_o = $signed(32'b00000000000000000000000000010110) <= $signed(n28566_o);
  /* rotator.vhdl:51:17  */
  assign n28571_o = n28568_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28572_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28573_o = {1'b0, n28572_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28575_o = $signed(32'b00000000000000000000000000010111) <= $signed(n28573_o);
  /* rotator.vhdl:51:17  */
  assign n28578_o = n28575_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28579_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28580_o = {1'b0, n28579_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28582_o = $signed(32'b00000000000000000000000000011000) <= $signed(n28580_o);
  /* rotator.vhdl:51:17  */
  assign n28585_o = n28582_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28586_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28587_o = {1'b0, n28586_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28589_o = $signed(32'b00000000000000000000000000011001) <= $signed(n28587_o);
  /* rotator.vhdl:51:17  */
  assign n28592_o = n28589_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28593_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28594_o = {1'b0, n28593_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28596_o = $signed(32'b00000000000000000000000000011010) <= $signed(n28594_o);
  /* rotator.vhdl:51:17  */
  assign n28599_o = n28596_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28600_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28601_o = {1'b0, n28600_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28603_o = $signed(32'b00000000000000000000000000011011) <= $signed(n28601_o);
  /* rotator.vhdl:51:17  */
  assign n28606_o = n28603_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28607_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28608_o = {1'b0, n28607_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28610_o = $signed(32'b00000000000000000000000000011100) <= $signed(n28608_o);
  /* rotator.vhdl:51:17  */
  assign n28613_o = n28610_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28614_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28615_o = {1'b0, n28614_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28617_o = $signed(32'b00000000000000000000000000011101) <= $signed(n28615_o);
  /* rotator.vhdl:51:17  */
  assign n28620_o = n28617_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28621_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28622_o = {1'b0, n28621_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28624_o = $signed(32'b00000000000000000000000000011110) <= $signed(n28622_o);
  /* rotator.vhdl:51:17  */
  assign n28627_o = n28624_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28628_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28629_o = {1'b0, n28628_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28631_o = $signed(32'b00000000000000000000000000011111) <= $signed(n28629_o);
  /* rotator.vhdl:51:17  */
  assign n28634_o = n28631_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28635_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28636_o = {1'b0, n28635_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28638_o = $signed(32'b00000000000000000000000000100000) <= $signed(n28636_o);
  /* rotator.vhdl:51:17  */
  assign n28641_o = n28638_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28642_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28643_o = {1'b0, n28642_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28645_o = $signed(32'b00000000000000000000000000100001) <= $signed(n28643_o);
  /* rotator.vhdl:51:17  */
  assign n28648_o = n28645_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28649_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28650_o = {1'b0, n28649_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28652_o = $signed(32'b00000000000000000000000000100010) <= $signed(n28650_o);
  /* rotator.vhdl:51:17  */
  assign n28655_o = n28652_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28656_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28657_o = {1'b0, n28656_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28659_o = $signed(32'b00000000000000000000000000100011) <= $signed(n28657_o);
  /* rotator.vhdl:51:17  */
  assign n28662_o = n28659_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28663_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28664_o = {1'b0, n28663_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28666_o = $signed(32'b00000000000000000000000000100100) <= $signed(n28664_o);
  /* rotator.vhdl:51:17  */
  assign n28669_o = n28666_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28670_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28671_o = {1'b0, n28670_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28673_o = $signed(32'b00000000000000000000000000100101) <= $signed(n28671_o);
  /* rotator.vhdl:51:17  */
  assign n28676_o = n28673_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28677_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28678_o = {1'b0, n28677_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28680_o = $signed(32'b00000000000000000000000000100110) <= $signed(n28678_o);
  /* rotator.vhdl:51:17  */
  assign n28683_o = n28680_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28684_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28685_o = {1'b0, n28684_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28687_o = $signed(32'b00000000000000000000000000100111) <= $signed(n28685_o);
  /* rotator.vhdl:51:17  */
  assign n28690_o = n28687_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28691_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28692_o = {1'b0, n28691_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28694_o = $signed(32'b00000000000000000000000000101000) <= $signed(n28692_o);
  /* rotator.vhdl:51:17  */
  assign n28697_o = n28694_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28698_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28699_o = {1'b0, n28698_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28701_o = $signed(32'b00000000000000000000000000101001) <= $signed(n28699_o);
  /* rotator.vhdl:51:17  */
  assign n28704_o = n28701_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28705_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28706_o = {1'b0, n28705_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28708_o = $signed(32'b00000000000000000000000000101010) <= $signed(n28706_o);
  /* rotator.vhdl:51:17  */
  assign n28711_o = n28708_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28712_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28713_o = {1'b0, n28712_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28715_o = $signed(32'b00000000000000000000000000101011) <= $signed(n28713_o);
  /* rotator.vhdl:51:17  */
  assign n28718_o = n28715_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28719_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28720_o = {1'b0, n28719_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28722_o = $signed(32'b00000000000000000000000000101100) <= $signed(n28720_o);
  /* rotator.vhdl:51:17  */
  assign n28725_o = n28722_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28726_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28727_o = {1'b0, n28726_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28729_o = $signed(32'b00000000000000000000000000101101) <= $signed(n28727_o);
  /* rotator.vhdl:51:17  */
  assign n28732_o = n28729_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28733_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28734_o = {1'b0, n28733_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28736_o = $signed(32'b00000000000000000000000000101110) <= $signed(n28734_o);
  /* rotator.vhdl:51:17  */
  assign n28739_o = n28736_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28740_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28741_o = {1'b0, n28740_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28743_o = $signed(32'b00000000000000000000000000101111) <= $signed(n28741_o);
  /* rotator.vhdl:51:17  */
  assign n28746_o = n28743_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28747_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28748_o = {1'b0, n28747_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28750_o = $signed(32'b00000000000000000000000000110000) <= $signed(n28748_o);
  /* rotator.vhdl:51:17  */
  assign n28753_o = n28750_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28754_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28755_o = {1'b0, n28754_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28757_o = $signed(32'b00000000000000000000000000110001) <= $signed(n28755_o);
  /* rotator.vhdl:51:17  */
  assign n28760_o = n28757_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28761_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28762_o = {1'b0, n28761_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28764_o = $signed(32'b00000000000000000000000000110010) <= $signed(n28762_o);
  /* rotator.vhdl:51:17  */
  assign n28767_o = n28764_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28768_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28769_o = {1'b0, n28768_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28771_o = $signed(32'b00000000000000000000000000110011) <= $signed(n28769_o);
  /* rotator.vhdl:51:17  */
  assign n28774_o = n28771_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28775_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28776_o = {1'b0, n28775_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28778_o = $signed(32'b00000000000000000000000000110100) <= $signed(n28776_o);
  /* rotator.vhdl:51:17  */
  assign n28781_o = n28778_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28782_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28783_o = {1'b0, n28782_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28785_o = $signed(32'b00000000000000000000000000110101) <= $signed(n28783_o);
  /* rotator.vhdl:51:17  */
  assign n28788_o = n28785_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28789_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28790_o = {1'b0, n28789_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28792_o = $signed(32'b00000000000000000000000000110110) <= $signed(n28790_o);
  /* rotator.vhdl:51:17  */
  assign n28795_o = n28792_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28796_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28797_o = {1'b0, n28796_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28799_o = $signed(32'b00000000000000000000000000110111) <= $signed(n28797_o);
  /* rotator.vhdl:51:17  */
  assign n28802_o = n28799_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28803_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28804_o = {1'b0, n28803_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28806_o = $signed(32'b00000000000000000000000000111000) <= $signed(n28804_o);
  /* rotator.vhdl:51:17  */
  assign n28809_o = n28806_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28810_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28811_o = {1'b0, n28810_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28813_o = $signed(32'b00000000000000000000000000111001) <= $signed(n28811_o);
  /* rotator.vhdl:51:17  */
  assign n28816_o = n28813_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28817_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28818_o = {1'b0, n28817_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28820_o = $signed(32'b00000000000000000000000000111010) <= $signed(n28818_o);
  /* rotator.vhdl:51:17  */
  assign n28823_o = n28820_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28824_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28825_o = {1'b0, n28824_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28827_o = $signed(32'b00000000000000000000000000111011) <= $signed(n28825_o);
  /* rotator.vhdl:51:17  */
  assign n28830_o = n28827_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28831_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28832_o = {1'b0, n28831_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28834_o = $signed(32'b00000000000000000000000000111100) <= $signed(n28832_o);
  /* rotator.vhdl:51:17  */
  assign n28837_o = n28834_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28838_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28839_o = {1'b0, n28838_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28841_o = $signed(32'b00000000000000000000000000111101) <= $signed(n28839_o);
  /* rotator.vhdl:51:17  */
  assign n28844_o = n28841_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28845_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28846_o = {1'b0, n28845_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28848_o = $signed(32'b00000000000000000000000000111110) <= $signed(n28846_o);
  /* rotator.vhdl:51:17  */
  assign n28851_o = n28848_o ? 1'b1 : 1'b0;
  /* rotator.vhdl:51:25  */
  assign n28852_o = {24'b0, me};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28853_o = {1'b0, n28852_o};  //  uext
  /* rotator.vhdl:51:22  */
  assign n28855_o = $signed(32'b00000000000000000000000000111111) <= $signed(n28853_o);
  /* rotator.vhdl:51:17  */
  assign n28858_o = n28855_o ? 1'b1 : 1'b0;
  assign n28859_o = {n28417_o, n28424_o, n28431_o, n28438_o, n28445_o, n28452_o, n28459_o, n28466_o, n28473_o, n28480_o, n28487_o, n28494_o, n28501_o, n28508_o, n28515_o, n28522_o, n28529_o, n28536_o, n28543_o, n28550_o, n28557_o, n28564_o, n28571_o, n28578_o, n28585_o, n28592_o, n28599_o, n28606_o, n28613_o, n28620_o, n28627_o, n28634_o, n28641_o, n28648_o, n28655_o, n28662_o, n28669_o, n28676_o, n28683_o, n28690_o, n28697_o, n28704_o, n28711_o, n28718_o, n28725_o, n28732_o, n28739_o, n28746_o, n28753_o, n28760_o, n28767_o, n28774_o, n28781_o, n28788_o, n28795_o, n28802_o, n28809_o, n28816_o, n28823_o, n28830_o, n28837_o, n28844_o, n28851_o, n28858_o};
  /* rotator.vhdl:49:9  */
  assign n28861_o = n28410_o ? n28859_o : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* rotator.vhdl:158:46  */
  assign n28863_o = ~clear_right;
  /* rotator.vhdl:158:30  */
  assign n28864_o = clear_left & n28863_o;
  /* rotator.vhdl:158:53  */
  assign n28865_o = n28864_o | right_shift;
  /* rotator.vhdl:160:47  */
  assign n28867_o = repl32[63];
  /* rotator.vhdl:160:37  */
  assign n28868_o = arith & n28867_o;
  /* rotator.vhdl:163:49  */
  assign n28870_o = mb[5:0];
  /* rotator.vhdl:163:76  */
  assign n28871_o = me[5:0];
  /* rotator.vhdl:163:63  */
  assign n28872_o = $unsigned(n28870_o) > $unsigned(n28871_o);
  /* rotator.vhdl:163:34  */
  assign n28873_o = clear_right & n28872_o;
  /* rotator.vhdl:163:13  */
  assign n28876_o = n28873_o ? 1'b1 : 1'b0;
  assign n28877_o = {1'b0, n28876_o};
  assign n28878_o = {1'b1, n28868_o};
  /* rotator.vhdl:158:9  */
  assign n28879_o = n28865_o ? n28878_o : n28877_o;
  /* rotator.vhdl:173:40  */
  assign n28880_o = mr & ml;
  /* rotator.vhdl:173:32  */
  assign n28881_o = rot & n28880_o;
  /* rotator.vhdl:173:68  */
  assign n28882_o = mr & ml;
  /* rotator.vhdl:173:60  */
  assign n28883_o = ~n28882_o;
  /* rotator.vhdl:173:56  */
  assign n28884_o = ra & n28883_o;
  /* rotator.vhdl:173:49  */
  assign n28885_o = n28881_o | n28884_o;
  /* rotator.vhdl:172:13  */
  assign n28887_o = output_mode == 2'b00;
  /* rotator.vhdl:175:40  */
  assign n28888_o = mr | ml;
  /* rotator.vhdl:175:32  */
  assign n28889_o = rot & n28888_o;
  /* rotator.vhdl:175:67  */
  assign n28890_o = mr | ml;
  /* rotator.vhdl:175:59  */
  assign n28891_o = ~n28890_o;
  /* rotator.vhdl:175:55  */
  assign n28892_o = ra & n28891_o;
  /* rotator.vhdl:175:48  */
  assign n28893_o = n28889_o | n28892_o;
  /* rotator.vhdl:174:13  */
  assign n28895_o = output_mode == 2'b01;
  /* rotator.vhdl:177:31  */
  assign n28896_o = rot & mr;
  /* rotator.vhdl:176:13  */
  assign n28898_o = output_mode == 2'b10;
  /* rotator.vhdl:179:34  */
  assign n28899_o = ~mr;
  /* rotator.vhdl:179:31  */
  assign n28900_o = rot | n28899_o;
  assign n28901_o = {n28898_o, n28895_o, n28887_o};
  /* rotator.vhdl:171:9  */
  always @*
    case (n28901_o)
      3'b100: n28902_o = n28896_o;
      3'b010: n28902_o = n28893_o;
      3'b001: n28902_o = n28885_o;
      default: n28902_o = n28900_o;
    endcase
  /* rotator.vhdl:183:24  */
  assign n28904_o = output_mode == 2'b11;
  /* rotator.vhdl:184:37  */
  assign n28905_o = ~ml;
  /* rotator.vhdl:184:33  */
  assign n28906_o = rs & n28905_o;
  /* rotator.vhdl:184:26  */
  assign n28907_o = |(n28906_o);
  /* rotator.vhdl:183:9  */
  assign n28909_o = n28904_o ? n28907_o : 1'b0;
endmodule

module control_3_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clk,
   input  rst,
   input  [1:0] complete_in_tag,
   input  complete_in_valid,
   input  valid_in,
   input  repeated,
   input  flush_in,
   input  busy_in,
   input  deferred,
   input  sgl_pipe_in,
   input  stop_mark_in,
   input  gpr_write_valid_in,
   input  [6:0] gpr_write_in,
   input  gpr_a_read_valid_in,
   input  [6:0] gpr_a_read_in,
   input  gpr_b_read_valid_in,
   input  [6:0] gpr_b_read_in,
   input  gpr_c_read_valid_in,
   input  [6:0] gpr_c_read_in,
   input  [1:0] execute_next_tag_tag,
   input  execute_next_tag_valid,
   input  [1:0] execute_next_cr_tag_tag,
   input  execute_next_cr_tag_valid,
   input  cr_read_in,
   input  cr_write_in,
   output valid_out,
   output stall_out,
   output stopped_out,
   output gpr_bypass_a,
   output gpr_bypass_b,
   output gpr_bypass_c,
   output cr_bypass,
   output [1:0] instr_tag_out_tag,
   output instr_tag_out_valid);
  wire [2:0] n26964_o;
  wire [2:0] n26965_o;
  wire [2:0] n26966_o;
  wire [1:0] n26975_o;
  wire n26976_o;
  reg [5:0] r_int;
  reg [5:0] rin_int;
  reg gpr_write_valid;
  reg cr_write_valid;
  wire [39:0] tag_regs;
  wire [2:0] instr_tag;
  wire gpr_tag_stall;
  wire cr_tag_stall;
  wire [1:0] curr_tag;
  wire [1:0] next_tag;
  wire [1:0] curr_cr_tag;
  wire n26983_o;
  wire n26986_o;
  wire [1:0] n26987_o;
  wire [31:0] n26988_o;
  wire n26990_o;
  wire n26991_o;
  wire n26994_o;
  wire n26995_o;
  wire n26996_o;
  wire n26997_o;
  wire [9:0] n26998_o;
  wire [6:0] n26999_o;
  wire n27000_o;
  wire n27001_o;
  wire n27008_o;
  wire n27009_o;
  wire n27010_o;
  wire [1:0] n27011_o;
  wire [31:0] n27012_o;
  wire n27014_o;
  wire n27015_o;
  wire [9:0] n27016_o;
  wire [6:0] n27017_o;
  wire [9:0] n27018_o;
  wire [9:0] n27019_o;
  wire n27020_o;
  wire n27021_o;
  wire [7:0] n27022_o;
  wire [7:0] n27023_o;
  wire [7:0] n27024_o;
  wire n27025_o;
  wire n27026_o;
  wire n27027_o;
  wire n27030_o;
  wire [1:0] n27031_o;
  wire [31:0] n27032_o;
  wire n27034_o;
  wire n27035_o;
  wire n27038_o;
  wire n27039_o;
  wire n27040_o;
  wire n27041_o;
  wire [9:0] n27042_o;
  wire [6:0] n27043_o;
  wire n27044_o;
  wire n27045_o;
  wire n27052_o;
  wire n27053_o;
  wire n27054_o;
  wire [1:0] n27055_o;
  wire [31:0] n27056_o;
  wire n27058_o;
  wire n27059_o;
  wire [9:0] n27060_o;
  wire [6:0] n27061_o;
  wire [9:0] n27062_o;
  wire [9:0] n27063_o;
  wire n27064_o;
  wire n27065_o;
  wire [7:0] n27066_o;
  wire [7:0] n27067_o;
  wire [7:0] n27068_o;
  wire n27069_o;
  wire n27070_o;
  wire n27071_o;
  wire n27074_o;
  wire [1:0] n27075_o;
  wire [31:0] n27076_o;
  wire n27078_o;
  wire n27079_o;
  wire n27082_o;
  wire n27083_o;
  wire n27084_o;
  wire n27085_o;
  wire [9:0] n27086_o;
  wire [6:0] n27087_o;
  wire n27088_o;
  wire n27089_o;
  wire n27096_o;
  wire n27097_o;
  wire n27098_o;
  wire [1:0] n27099_o;
  wire [31:0] n27100_o;
  wire n27102_o;
  wire n27103_o;
  wire [9:0] n27104_o;
  wire [6:0] n27105_o;
  wire [9:0] n27106_o;
  wire [9:0] n27107_o;
  wire n27108_o;
  wire n27109_o;
  wire [7:0] n27110_o;
  wire [7:0] n27111_o;
  wire [7:0] n27112_o;
  wire n27113_o;
  wire n27114_o;
  wire n27115_o;
  wire n27118_o;
  wire [1:0] n27119_o;
  wire [31:0] n27120_o;
  wire n27122_o;
  wire n27123_o;
  wire n27126_o;
  wire n27127_o;
  wire n27128_o;
  wire n27129_o;
  wire [9:0] n27130_o;
  wire [6:0] n27131_o;
  wire n27132_o;
  wire n27133_o;
  wire n27140_o;
  wire n27141_o;
  wire n27142_o;
  wire [1:0] n27143_o;
  wire [31:0] n27144_o;
  wire n27146_o;
  wire n27147_o;
  wire [9:0] n27148_o;
  wire [6:0] n27149_o;
  wire [9:0] n27150_o;
  wire [9:0] n27151_o;
  wire n27152_o;
  wire n27153_o;
  wire [7:0] n27154_o;
  wire [7:0] n27155_o;
  wire [7:0] n27156_o;
  wire n27157_o;
  wire n27158_o;
  wire [1:0] n27159_o;
  wire [1:0] n27160_o;
  wire [1:0] n27162_o;
  wire [1:0] n27164_o;
  wire [39:0] n27166_o;
  wire [9:0] n27184_o;
  wire n27185_o;
  wire [9:0] n27186_o;
  wire n27187_o;
  wire n27188_o;
  wire [9:0] n27189_o;
  wire [6:0] n27190_o;
  wire n27191_o;
  wire n27192_o;
  wire [2:0] n27194_o;
  localparam [2:0] n27195_o = 3'b000;
  wire [2:0] n27196_o;
  wire [9:0] n27198_o;
  wire n27199_o;
  wire [9:0] n27200_o;
  wire n27201_o;
  wire n27202_o;
  wire [9:0] n27203_o;
  wire [6:0] n27204_o;
  wire n27205_o;
  wire n27206_o;
  wire [2:0] n27208_o;
  wire [2:0] n27209_o;
  wire [9:0] n27210_o;
  wire n27211_o;
  wire [9:0] n27212_o;
  wire n27213_o;
  wire n27214_o;
  wire [9:0] n27215_o;
  wire [6:0] n27216_o;
  wire n27217_o;
  wire n27218_o;
  wire [2:0] n27220_o;
  wire [2:0] n27221_o;
  wire [9:0] n27222_o;
  wire n27223_o;
  wire [9:0] n27224_o;
  wire n27225_o;
  wire n27226_o;
  wire [9:0] n27227_o;
  wire [6:0] n27228_o;
  wire n27229_o;
  wire n27230_o;
  wire [2:0] n27232_o;
  wire [2:0] n27233_o;
  wire n27239_o;
  wire n27240_o;
  wire n27241_o;
  wire [1:0] n27242_o;
  wire [31:0] n27243_o;
  wire [1:0] n27244_o;
  wire [31:0] n27245_o;
  wire n27246_o;
  wire n27247_o;
  wire n27249_o;
  wire n27250_o;
  wire n27251_o;
  wire n27252_o;
  wire n27253_o;
  wire n27254_o;
  wire n27255_o;
  wire n27256_o;
  wire n27257_o;
  wire n27258_o;
  wire [1:0] n27259_o;
  wire [1:0] n27260_o;
  wire [1:0] n27261_o;
  wire [1:0] n27262_o;
  wire [1:0] n27263_o;
  wire [1:0] n27264_o;
  wire [1:0] n27265_o;
  wire [1:0] n27266_o;
  wire [1:0] n27267_o;
  wire [9:0] n27268_o;
  wire n27269_o;
  wire [9:0] n27270_o;
  wire n27271_o;
  wire n27272_o;
  wire [9:0] n27273_o;
  wire [6:0] n27274_o;
  wire n27275_o;
  wire n27276_o;
  wire [2:0] n27278_o;
  localparam [2:0] n27279_o = 3'b000;
  wire [2:0] n27280_o;
  wire [9:0] n27282_o;
  wire n27283_o;
  wire [9:0] n27284_o;
  wire n27285_o;
  wire n27286_o;
  wire [9:0] n27287_o;
  wire [6:0] n27288_o;
  wire n27289_o;
  wire n27290_o;
  wire [2:0] n27292_o;
  wire [2:0] n27293_o;
  wire [9:0] n27294_o;
  wire n27295_o;
  wire [9:0] n27296_o;
  wire n27297_o;
  wire n27298_o;
  wire [9:0] n27299_o;
  wire [6:0] n27300_o;
  wire n27301_o;
  wire n27302_o;
  wire [2:0] n27304_o;
  wire [2:0] n27305_o;
  wire [9:0] n27306_o;
  wire n27307_o;
  wire [9:0] n27308_o;
  wire n27309_o;
  wire n27310_o;
  wire [9:0] n27311_o;
  wire [6:0] n27312_o;
  wire n27313_o;
  wire n27314_o;
  wire [2:0] n27316_o;
  wire [2:0] n27317_o;
  wire n27323_o;
  wire n27324_o;
  wire n27325_o;
  wire [1:0] n27326_o;
  wire [31:0] n27327_o;
  wire [1:0] n27328_o;
  wire [31:0] n27329_o;
  wire n27330_o;
  wire n27331_o;
  wire n27333_o;
  wire n27334_o;
  wire n27335_o;
  wire n27336_o;
  wire n27337_o;
  wire n27338_o;
  wire n27339_o;
  wire n27340_o;
  wire n27341_o;
  wire n27342_o;
  wire [1:0] n27343_o;
  wire [1:0] n27344_o;
  wire [1:0] n27345_o;
  wire [1:0] n27346_o;
  wire [1:0] n27347_o;
  wire [1:0] n27348_o;
  wire [1:0] n27349_o;
  wire [1:0] n27350_o;
  wire [1:0] n27351_o;
  wire [9:0] n27352_o;
  wire n27353_o;
  wire [9:0] n27354_o;
  wire n27355_o;
  wire n27356_o;
  wire [9:0] n27357_o;
  wire [6:0] n27358_o;
  wire n27359_o;
  wire n27360_o;
  wire [2:0] n27362_o;
  localparam [2:0] n27363_o = 3'b000;
  wire [2:0] n27364_o;
  wire [9:0] n27366_o;
  wire n27367_o;
  wire [9:0] n27368_o;
  wire n27369_o;
  wire n27370_o;
  wire [9:0] n27371_o;
  wire [6:0] n27372_o;
  wire n27373_o;
  wire n27374_o;
  wire [2:0] n27376_o;
  wire [2:0] n27377_o;
  wire [9:0] n27378_o;
  wire n27379_o;
  wire [9:0] n27380_o;
  wire n27381_o;
  wire n27382_o;
  wire [9:0] n27383_o;
  wire [6:0] n27384_o;
  wire n27385_o;
  wire n27386_o;
  wire [2:0] n27388_o;
  wire [2:0] n27389_o;
  wire [9:0] n27390_o;
  wire n27391_o;
  wire [9:0] n27392_o;
  wire n27393_o;
  wire n27394_o;
  wire [9:0] n27395_o;
  wire [6:0] n27396_o;
  wire n27397_o;
  wire n27398_o;
  wire [2:0] n27400_o;
  wire [2:0] n27401_o;
  wire n27407_o;
  wire n27408_o;
  wire n27409_o;
  wire [1:0] n27410_o;
  wire [31:0] n27411_o;
  wire [1:0] n27412_o;
  wire [31:0] n27413_o;
  wire n27414_o;
  wire n27415_o;
  wire n27417_o;
  wire n27418_o;
  wire n27419_o;
  wire n27420_o;
  wire n27421_o;
  wire n27422_o;
  wire n27423_o;
  wire n27424_o;
  wire n27425_o;
  wire n27426_o;
  wire [1:0] n27427_o;
  wire [1:0] n27428_o;
  wire [1:0] n27429_o;
  wire [1:0] n27430_o;
  wire [1:0] n27431_o;
  wire [1:0] n27432_o;
  wire [1:0] n27433_o;
  wire [1:0] n27434_o;
  wire [1:0] n27435_o;
  wire n27441_o;
  wire [2:0] n27442_o;
  wire n27443_o;
  wire n27444_o;
  wire [1:0] n27445_o;
  wire [31:0] n27446_o;
  wire [2:0] n27447_o;
  wire [1:0] n27448_o;
  wire [31:0] n27449_o;
  wire n27450_o;
  wire n27451_o;
  wire n27453_o;
  wire n27456_o;
  wire n27463_o;
  wire [2:0] n27464_o;
  wire n27465_o;
  wire n27466_o;
  wire [1:0] n27467_o;
  wire [31:0] n27468_o;
  wire [2:0] n27469_o;
  wire [1:0] n27470_o;
  wire [31:0] n27471_o;
  wire n27472_o;
  wire n27473_o;
  wire n27475_o;
  wire n27478_o;
  wire n27485_o;
  wire [2:0] n27486_o;
  wire n27487_o;
  wire n27488_o;
  wire [1:0] n27489_o;
  wire [31:0] n27490_o;
  wire [2:0] n27491_o;
  wire [1:0] n27492_o;
  wire [31:0] n27493_o;
  wire n27494_o;
  wire n27495_o;
  wire n27497_o;
  wire n27500_o;
  wire [2:0] n27502_o;
  wire n27503_o;
  wire n27504_o;
  wire n27505_o;
  wire [2:0] n27506_o;
  wire n27507_o;
  wire n27508_o;
  wire n27509_o;
  wire n27510_o;
  wire [2:0] n27511_o;
  wire n27512_o;
  wire n27513_o;
  wire n27514_o;
  wire n27515_o;
  wire n27516_o;
  wire n27517_o;
  wire n27518_o;
  wire [31:0] n27519_o;
  wire [31:0] n27521_o;
  wire [1:0] n27522_o;
  wire [1:0] n27524_o;
  wire [1:0] n27526_o;
  wire n27529_o;
  wire n27530_o;
  wire [2:0] n27536_o;
  wire n27537_o;
  wire n27538_o;
  wire n27539_o;
  wire [2:0] n27540_o;
  wire [1:0] n27541_o;
  wire [31:0] n27542_o;
  wire [1:0] n27543_o;
  wire [31:0] n27544_o;
  wire n27545_o;
  wire n27546_o;
  wire n27548_o;
  wire n27554_o;
  wire [2:0] n27555_o;
  wire n27556_o;
  wire n27557_o;
  wire [1:0] n27558_o;
  wire [31:0] n27559_o;
  wire [2:0] n27560_o;
  wire [1:0] n27561_o;
  wire [31:0] n27562_o;
  wire n27563_o;
  wire n27564_o;
  wire n27566_o;
  wire n27569_o;
  wire [2:0] n27571_o;
  wire n27572_o;
  wire n27573_o;
  wire n27574_o;
  wire n27589_o;
  wire n27590_o;
  wire n27592_o;
  wire [3:0] n27593_o;
  wire [31:0] n27594_o;
  wire [31:0] n27596_o;
  wire [3:0] n27597_o;
  wire [3:0] n27598_o;
  wire [3:0] n27599_o;
  wire [3:0] n27600_o;
  wire [1:0] n27601_o;
  wire [3:0] n27602_o;
  wire [31:0] n27603_o;
  wire n27605_o;
  wire n27607_o;
  wire n27610_o;
  localparam [5:0] n27612_o = 6'b000000;
  wire [5:0] n27613_o;
  wire [5:0] n27614_o;
  wire n27616_o;
  wire [3:0] n27617_o;
  wire [31:0] n27618_o;
  wire n27620_o;
  wire n27621_o;
  wire n27624_o;
  wire [1:0] n27626_o;
  wire [3:0] n27627_o;
  wire [31:0] n27628_o;
  wire n27630_o;
  wire [1:0] n27633_o;
  wire n27635_o;
  wire n27636_o;
  wire [1:0] n27637_o;
  wire [1:0] n27638_o;
  wire [1:0] n27639_o;
  wire [1:0] n27640_o;
  wire n27641_o;
  wire [1:0] n27642_o;
  wire [1:0] n27643_o;
  wire [1:0] n27644_o;
  wire [1:0] n27645_o;
  wire n27646_o;
  wire n27648_o;
  wire [3:0] n27649_o;
  wire [31:0] n27650_o;
  wire n27652_o;
  wire [1:0] n27654_o;
  wire [1:0] n27655_o;
  wire [1:0] n27656_o;
  wire [1:0] n27657_o;
  wire n27659_o;
  wire n27661_o;
  wire [3:0] n27662_o;
  wire [31:0] n27663_o;
  wire n27665_o;
  wire [3:0] n27667_o;
  wire [3:0] n27668_o;
  wire [3:0] n27669_o;
  wire [5:0] n27670_o;
  wire [3:0] n27671_o;
  wire [31:0] n27672_o;
  wire n27674_o;
  wire [1:0] n27677_o;
  wire n27679_o;
  wire n27680_o;
  wire [1:0] n27681_o;
  wire n27682_o;
  wire n27683_o;
  wire n27684_o;
  wire [1:0] n27685_o;
  wire [1:0] n27686_o;
  wire [1:0] n27687_o;
  wire [1:0] n27688_o;
  wire n27690_o;
  wire n27692_o;
  wire [2:0] n27693_o;
  reg [1:0] n27695_o;
  wire [3:0] n27696_o;
  wire [3:0] n27697_o;
  wire [3:0] n27698_o;
  reg n27700_o;
  wire n27702_o;
  wire n27703_o;
  wire n27704_o;
  wire n27705_o;
  wire n27706_o;
  wire [5:0] n27707_o;
  wire [3:0] n27708_o;
  wire [31:0] n27709_o;
  wire [31:0] n27711_o;
  wire [3:0] n27712_o;
  wire [3:0] n27713_o;
  wire n27714_o;
  wire [5:0] n27715_o;
  reg [5:0] n27719_q;
  reg [39:0] n27720_q;
  wire [2:0] n27721_o;
  reg [1:0] n27722_q;
  reg [1:0] n27723_q;
  wire [9:0] n27724_o;
  wire [9:0] n27725_o;
  wire [9:0] n27726_o;
  wire [9:0] n27727_o;
  wire [1:0] n27728_o;
  reg [9:0] n27729_o;
  assign valid_out = n27702_o;
  assign stall_out = n27714_o;
  assign stopped_out = n27624_o;
  assign gpr_bypass_a = n27456_o;
  assign gpr_bypass_b = n27478_o;
  assign gpr_bypass_c = n27500_o;
  assign cr_bypass = n27569_o;
  assign instr_tag_out_tag = n26975_o;
  assign instr_tag_out_valid = n26976_o;
  /* asic/cache_ram.vhdl:19:9  */
  assign n26964_o = {complete_in_valid, complete_in_tag};
  /* spi_rxtx.vhdl:154:14  */
  assign n26965_o = {execute_next_tag_valid, execute_next_tag_tag};
  /* asic/cache_ram.vhdl:75:9  */
  assign n26966_o = {execute_next_cr_tag_valid, execute_next_cr_tag_tag};
  /* spi_rxtx.vhdl:150:14  */
  assign n26975_o = instr_tag[1:0];
  assign n26976_o = instr_tag[2];
  /* control.vhdl:65:12  */
  always @*
    r_int = n27719_q; // (isignal)
  initial
    r_int = 6'b000000;
  /* control.vhdl:65:19  */
  always @*
    rin_int = n27715_o; // (isignal)
  initial
    rin_int = 6'b000000;
  /* control.vhdl:67:12  */
  always @*
    gpr_write_valid = n27703_o; // (isignal)
  initial
    gpr_write_valid = 1'b0;
  /* control.vhdl:68:12  */
  always @*
    cr_write_valid = n27704_o; // (isignal)
  initial
    cr_write_valid = 1'b0;
  /* control.vhdl:78:12  */
  assign tag_regs = n27720_q; // (signal)
  /* control.vhdl:80:12  */
  assign instr_tag = n27721_o; // (signal)
  /* control.vhdl:82:12  */
  assign gpr_tag_stall = n27515_o; // (signal)
  /* control.vhdl:83:12  */
  assign cr_tag_stall = n27574_o; // (signal)
  /* control.vhdl:85:12  */
  assign curr_tag = n27722_q; // (signal)
  /* control.vhdl:86:12  */
  assign next_tag = n27524_o; // (signal)
  /* control.vhdl:88:12  */
  assign curr_cr_tag = n27723_q; // (signal)
  /* control.vhdl:98:30  */
  assign n26983_o = rst | flush_in;
  /* control.vhdl:102:36  */
  assign n26986_o = n26964_o[2];
  /* control.vhdl:102:68  */
  assign n26987_o = n26964_o[1:0];
  /* control.vhdl:102:54  */
  assign n26988_o = {30'b0, n26987_o};  //  uext
  /* control.vhdl:102:54  */
  assign n26990_o = 32'b00000000000000000000000000000000 == n26988_o;
  /* control.vhdl:102:48  */
  assign n26991_o = n26986_o & n26990_o;
  /* spi_rxtx.vhdl:146:14  */
  assign n26994_o = tag_regs[30];
  /* control.vhdl:102:21  */
  assign n26995_o = n26991_o ? 1'b0 : n26994_o;
  /* spi_rxtx.vhdl:146:14  */
  assign n26996_o = tag_regs[39];
  /* control.vhdl:102:21  */
  assign n26997_o = n26991_o ? 1'b0 : n26996_o;
  /* control.vhdl:107:58  */
  assign n26998_o = tag_regs[39:30];
  /* control.vhdl:107:62  */
  assign n26999_o = n26998_o[7:1];
  /* control.vhdl:107:66  */
  assign n27000_o = n26999_o == gpr_write_in;
  /* control.vhdl:107:46  */
  assign n27001_o = gpr_write_valid & n27000_o;
  assign n27008_o = tag_regs[38];
  /* control.vhdl:107:21  */
  assign n27009_o = n27001_o ? 1'b0 : n27008_o;
  /* control.vhdl:113:34  */
  assign n27010_o = instr_tag[2];
  /* control.vhdl:113:64  */
  assign n27011_o = instr_tag[1:0];
  /* control.vhdl:113:52  */
  assign n27012_o = {30'b0, n27011_o};  //  uext
  /* control.vhdl:113:52  */
  assign n27014_o = 32'b00000000000000000000000000000000 == n27012_o;
  /* control.vhdl:113:46  */
  assign n27015_o = n27010_o & n27014_o;
  assign n27016_o = {cr_write_valid, gpr_write_valid, gpr_write_in, gpr_write_valid};
  assign n27017_o = tag_regs[37:31];
  assign n27018_o = {n26997_o, n27009_o, n27017_o, n26995_o};
  /* control.vhdl:113:21  */
  assign n27019_o = n27015_o ? n27016_o : n27018_o;
  assign n27020_o = n27019_o[0];
  /* control.vhdl:98:17  */
  assign n27021_o = n26983_o ? 1'b0 : n27020_o;
  assign n27022_o = n27019_o[8:1];
  assign n27023_o = tag_regs[38:31];
  /* control.vhdl:98:17  */
  assign n27024_o = n26983_o ? n27023_o : n27022_o;
  assign n27025_o = n27019_o[9];
  /* control.vhdl:98:17  */
  assign n27026_o = n26983_o ? 1'b0 : n27025_o;
  /* control.vhdl:98:30  */
  assign n27027_o = rst | flush_in;
  /* control.vhdl:102:36  */
  assign n27030_o = n26964_o[2];
  /* control.vhdl:102:68  */
  assign n27031_o = n26964_o[1:0];
  /* control.vhdl:102:54  */
  assign n27032_o = {30'b0, n27031_o};  //  uext
  /* control.vhdl:102:54  */
  assign n27034_o = 32'b00000000000000000000000000000001 == n27032_o;
  /* control.vhdl:102:48  */
  assign n27035_o = n27030_o & n27034_o;
  assign n27038_o = tag_regs[20];
  /* control.vhdl:102:21  */
  assign n27039_o = n27035_o ? 1'b0 : n27038_o;
  assign n27040_o = tag_regs[29];
  /* control.vhdl:102:21  */
  assign n27041_o = n27035_o ? 1'b0 : n27040_o;
  /* control.vhdl:107:58  */
  assign n27042_o = tag_regs[29:20];
  /* control.vhdl:107:62  */
  assign n27043_o = n27042_o[7:1];
  /* control.vhdl:107:66  */
  assign n27044_o = n27043_o == gpr_write_in;
  /* control.vhdl:107:46  */
  assign n27045_o = gpr_write_valid & n27044_o;
  assign n27052_o = tag_regs[28];
  /* control.vhdl:107:21  */
  assign n27053_o = n27045_o ? 1'b0 : n27052_o;
  /* control.vhdl:113:34  */
  assign n27054_o = instr_tag[2];
  /* control.vhdl:113:64  */
  assign n27055_o = instr_tag[1:0];
  /* control.vhdl:113:52  */
  assign n27056_o = {30'b0, n27055_o};  //  uext
  /* control.vhdl:113:52  */
  assign n27058_o = 32'b00000000000000000000000000000001 == n27056_o;
  /* control.vhdl:113:46  */
  assign n27059_o = n27054_o & n27058_o;
  assign n27060_o = {cr_write_valid, gpr_write_valid, gpr_write_in, gpr_write_valid};
  assign n27061_o = tag_regs[27:21];
  assign n27062_o = {n27041_o, n27053_o, n27061_o, n27039_o};
  /* control.vhdl:113:21  */
  assign n27063_o = n27059_o ? n27060_o : n27062_o;
  assign n27064_o = n27063_o[0];
  /* control.vhdl:98:17  */
  assign n27065_o = n27027_o ? 1'b0 : n27064_o;
  assign n27066_o = n27063_o[8:1];
  assign n27067_o = tag_regs[28:21];
  /* control.vhdl:98:17  */
  assign n27068_o = n27027_o ? n27067_o : n27066_o;
  assign n27069_o = n27063_o[9];
  /* control.vhdl:98:17  */
  assign n27070_o = n27027_o ? 1'b0 : n27069_o;
  /* control.vhdl:98:30  */
  assign n27071_o = rst | flush_in;
  /* control.vhdl:102:36  */
  assign n27074_o = n26964_o[2];
  /* control.vhdl:102:68  */
  assign n27075_o = n26964_o[1:0];
  /* control.vhdl:102:54  */
  assign n27076_o = {30'b0, n27075_o};  //  uext
  /* control.vhdl:102:54  */
  assign n27078_o = 32'b00000000000000000000000000000010 == n27076_o;
  /* control.vhdl:102:48  */
  assign n27079_o = n27074_o & n27078_o;
  assign n27082_o = tag_regs[10];
  /* control.vhdl:102:21  */
  assign n27083_o = n27079_o ? 1'b0 : n27082_o;
  assign n27084_o = tag_regs[19];
  /* control.vhdl:102:21  */
  assign n27085_o = n27079_o ? 1'b0 : n27084_o;
  /* control.vhdl:107:58  */
  assign n27086_o = tag_regs[19:10];
  /* control.vhdl:107:62  */
  assign n27087_o = n27086_o[7:1];
  /* control.vhdl:107:66  */
  assign n27088_o = n27087_o == gpr_write_in;
  /* control.vhdl:107:46  */
  assign n27089_o = gpr_write_valid & n27088_o;
  assign n27096_o = tag_regs[18];
  /* control.vhdl:107:21  */
  assign n27097_o = n27089_o ? 1'b0 : n27096_o;
  /* control.vhdl:113:34  */
  assign n27098_o = instr_tag[2];
  /* control.vhdl:113:64  */
  assign n27099_o = instr_tag[1:0];
  /* control.vhdl:113:52  */
  assign n27100_o = {30'b0, n27099_o};  //  uext
  /* control.vhdl:113:52  */
  assign n27102_o = 32'b00000000000000000000000000000010 == n27100_o;
  /* control.vhdl:113:46  */
  assign n27103_o = n27098_o & n27102_o;
  assign n27104_o = {cr_write_valid, gpr_write_valid, gpr_write_in, gpr_write_valid};
  assign n27105_o = tag_regs[17:11];
  assign n27106_o = {n27085_o, n27097_o, n27105_o, n27083_o};
  /* control.vhdl:113:21  */
  assign n27107_o = n27103_o ? n27104_o : n27106_o;
  assign n27108_o = n27107_o[0];
  /* control.vhdl:98:17  */
  assign n27109_o = n27071_o ? 1'b0 : n27108_o;
  assign n27110_o = n27107_o[8:1];
  assign n27111_o = tag_regs[18:11];
  /* control.vhdl:98:17  */
  assign n27112_o = n27071_o ? n27111_o : n27110_o;
  assign n27113_o = n27107_o[9];
  /* control.vhdl:98:17  */
  assign n27114_o = n27071_o ? 1'b0 : n27113_o;
  /* control.vhdl:98:30  */
  assign n27115_o = rst | flush_in;
  /* control.vhdl:102:36  */
  assign n27118_o = n26964_o[2];
  /* control.vhdl:102:68  */
  assign n27119_o = n26964_o[1:0];
  /* control.vhdl:102:54  */
  assign n27120_o = {30'b0, n27119_o};  //  uext
  /* control.vhdl:102:54  */
  assign n27122_o = 32'b00000000000000000000000000000011 == n27120_o;
  /* control.vhdl:102:48  */
  assign n27123_o = n27118_o & n27122_o;
  assign n27126_o = tag_regs[0];
  /* control.vhdl:102:21  */
  assign n27127_o = n27123_o ? 1'b0 : n27126_o;
  assign n27128_o = tag_regs[9];
  /* control.vhdl:102:21  */
  assign n27129_o = n27123_o ? 1'b0 : n27128_o;
  /* control.vhdl:107:58  */
  assign n27130_o = tag_regs[9:0];
  /* control.vhdl:107:62  */
  assign n27131_o = n27130_o[7:1];
  /* control.vhdl:107:66  */
  assign n27132_o = n27131_o == gpr_write_in;
  /* control.vhdl:107:46  */
  assign n27133_o = gpr_write_valid & n27132_o;
  assign n27140_o = tag_regs[8];
  /* control.vhdl:107:21  */
  assign n27141_o = n27133_o ? 1'b0 : n27140_o;
  /* control.vhdl:113:34  */
  assign n27142_o = instr_tag[2];
  /* control.vhdl:113:64  */
  assign n27143_o = instr_tag[1:0];
  /* control.vhdl:113:52  */
  assign n27144_o = {30'b0, n27143_o};  //  uext
  /* control.vhdl:113:52  */
  assign n27146_o = 32'b00000000000000000000000000000011 == n27144_o;
  /* control.vhdl:113:46  */
  assign n27147_o = n27142_o & n27146_o;
  assign n27148_o = {cr_write_valid, gpr_write_valid, gpr_write_in, gpr_write_valid};
  assign n27149_o = tag_regs[7:1];
  assign n27150_o = {n27129_o, n27141_o, n27149_o, n27127_o};
  /* control.vhdl:113:21  */
  assign n27151_o = n27147_o ? n27148_o : n27150_o;
  assign n27152_o = n27151_o[0];
  /* control.vhdl:98:17  */
  assign n27153_o = n27115_o ? 1'b0 : n27152_o;
  assign n27154_o = n27151_o[8:1];
  assign n27155_o = tag_regs[8:1];
  /* control.vhdl:98:17  */
  assign n27156_o = n27115_o ? n27155_o : n27154_o;
  assign n27157_o = n27151_o[9];
  /* control.vhdl:98:17  */
  assign n27158_o = n27115_o ? 1'b0 : n27157_o;
  /* control.vhdl:130:46  */
  assign n27159_o = instr_tag[1:0];
  /* control.vhdl:129:17  */
  assign n27160_o = cr_write_valid ? n27159_o : curr_cr_tag;
  /* control.vhdl:124:13  */
  assign n27162_o = rst ? 2'b00 : next_tag;
  /* control.vhdl:124:13  */
  assign n27164_o = rst ? 2'b00 : n27160_o;
  assign n27166_o = {n27026_o, n27024_o, n27021_o, n27070_o, n27068_o, n27065_o, n27114_o, n27112_o, n27109_o, n27158_o, n27156_o, n27153_o};
  /* control.vhdl:152:24  */
  assign n27184_o = tag_regs[39:30];
  /* control.vhdl:152:28  */
  assign n27185_o = n27184_o[0];
  /* control.vhdl:152:53  */
  assign n27186_o = tag_regs[39:30];
  /* control.vhdl:152:57  */
  assign n27187_o = n27186_o[8];
  /* control.vhdl:152:41  */
  assign n27188_o = n27185_o & n27187_o;
  /* control.vhdl:152:82  */
  assign n27189_o = tag_regs[39:30];
  /* control.vhdl:152:86  */
  assign n27190_o = n27189_o[7:1];
  /* control.vhdl:152:90  */
  assign n27191_o = n27190_o == gpr_a_read_in;
  /* control.vhdl:152:70  */
  assign n27192_o = n27188_o & n27191_o;
  assign n27194_o = {gpr_a_read_valid_in, 2'b00};
  /* control.vhdl:152:13  */
  assign n27196_o = n27192_o ? n27194_o : 3'b000;
  /* control.vhdl:152:24  */
  assign n27198_o = tag_regs[29:20];
  /* control.vhdl:152:28  */
  assign n27199_o = n27198_o[0];
  /* control.vhdl:152:53  */
  assign n27200_o = tag_regs[29:20];
  /* control.vhdl:152:57  */
  assign n27201_o = n27200_o[8];
  /* control.vhdl:152:41  */
  assign n27202_o = n27199_o & n27201_o;
  /* control.vhdl:152:82  */
  assign n27203_o = tag_regs[29:20];
  /* control.vhdl:152:86  */
  assign n27204_o = n27203_o[7:1];
  /* control.vhdl:152:90  */
  assign n27205_o = n27204_o == gpr_a_read_in;
  /* control.vhdl:152:70  */
  assign n27206_o = n27202_o & n27205_o;
  assign n27208_o = {gpr_a_read_valid_in, 2'b01};
  /* control.vhdl:152:13  */
  assign n27209_o = n27206_o ? n27208_o : n27196_o;
  /* control.vhdl:152:24  */
  assign n27210_o = tag_regs[19:10];
  /* control.vhdl:152:28  */
  assign n27211_o = n27210_o[0];
  /* control.vhdl:152:53  */
  assign n27212_o = tag_regs[19:10];
  /* control.vhdl:152:57  */
  assign n27213_o = n27212_o[8];
  /* control.vhdl:152:41  */
  assign n27214_o = n27211_o & n27213_o;
  /* control.vhdl:152:82  */
  assign n27215_o = tag_regs[19:10];
  /* control.vhdl:152:86  */
  assign n27216_o = n27215_o[7:1];
  /* control.vhdl:152:90  */
  assign n27217_o = n27216_o == gpr_a_read_in;
  /* control.vhdl:152:70  */
  assign n27218_o = n27214_o & n27217_o;
  assign n27220_o = {gpr_a_read_valid_in, 2'b10};
  /* control.vhdl:152:13  */
  assign n27221_o = n27218_o ? n27220_o : n27209_o;
  /* control.vhdl:152:24  */
  assign n27222_o = tag_regs[9:0];
  /* control.vhdl:152:28  */
  assign n27223_o = n27222_o[0];
  /* control.vhdl:152:53  */
  assign n27224_o = tag_regs[9:0];
  /* control.vhdl:152:57  */
  assign n27225_o = n27224_o[8];
  /* control.vhdl:152:41  */
  assign n27226_o = n27223_o & n27225_o;
  /* control.vhdl:152:82  */
  assign n27227_o = tag_regs[9:0];
  /* control.vhdl:152:86  */
  assign n27228_o = n27227_o[7:1];
  /* control.vhdl:152:90  */
  assign n27229_o = n27228_o == gpr_a_read_in;
  /* control.vhdl:152:70  */
  assign n27230_o = n27226_o & n27229_o;
  assign n27232_o = {gpr_a_read_valid_in, 2'b11};
  /* control.vhdl:152:13  */
  assign n27233_o = n27230_o ? n27232_o : n27221_o;
  /* common.vhdl:785:21  */
  assign n27239_o = n27233_o[2];
  /* common.vhdl:785:42  */
  assign n27240_o = n26964_o[2];
  /* common.vhdl:785:33  */
  assign n27241_o = n27239_o & n27240_o;
  /* common.vhdl:785:63  */
  assign n27242_o = n27233_o[1:0];
  /* common.vhdl:785:67  */
  assign n27243_o = {30'b0, n27242_o};  //  uext
  /* common.vhdl:785:74  */
  assign n27244_o = n26964_o[1:0];
  /* common.vhdl:785:67  */
  assign n27245_o = {30'b0, n27244_o};  //  uext
  /* common.vhdl:785:67  */
  assign n27246_o = n27243_o == n27245_o;
  /* common.vhdl:785:54  */
  assign n27247_o = n27241_o & n27246_o;
  assign n27249_o = n27232_o[2];
  assign n27250_o = n27220_o[2];
  assign n27251_o = n27208_o[2];
  assign n27252_o = n27194_o[2];
  assign n27253_o = n27195_o[2];
  /* control.vhdl:152:13  */
  assign n27254_o = n27192_o ? n27252_o : n27253_o;
  /* control.vhdl:152:13  */
  assign n27255_o = n27206_o ? n27251_o : n27254_o;
  /* control.vhdl:152:13  */
  assign n27256_o = n27218_o ? n27250_o : n27255_o;
  /* control.vhdl:152:13  */
  assign n27257_o = n27230_o ? n27249_o : n27256_o;
  /* control.vhdl:157:9  */
  assign n27258_o = n27247_o ? 1'b0 : n27257_o;
  assign n27259_o = n27232_o[1:0];
  assign n27260_o = n27220_o[1:0];
  assign n27261_o = n27208_o[1:0];
  assign n27262_o = n27194_o[1:0];
  assign n27263_o = n27195_o[1:0];
  /* control.vhdl:152:13  */
  assign n27264_o = n27192_o ? n27262_o : n27263_o;
  /* control.vhdl:152:13  */
  assign n27265_o = n27206_o ? n27261_o : n27264_o;
  /* control.vhdl:152:13  */
  assign n27266_o = n27218_o ? n27260_o : n27265_o;
  /* control.vhdl:152:13  */
  assign n27267_o = n27230_o ? n27259_o : n27266_o;
  /* control.vhdl:162:24  */
  assign n27268_o = tag_regs[39:30];
  /* control.vhdl:162:28  */
  assign n27269_o = n27268_o[0];
  /* control.vhdl:162:53  */
  assign n27270_o = tag_regs[39:30];
  /* control.vhdl:162:57  */
  assign n27271_o = n27270_o[8];
  /* control.vhdl:162:41  */
  assign n27272_o = n27269_o & n27271_o;
  /* control.vhdl:162:82  */
  assign n27273_o = tag_regs[39:30];
  /* control.vhdl:162:86  */
  assign n27274_o = n27273_o[7:1];
  /* control.vhdl:162:90  */
  assign n27275_o = n27274_o == gpr_b_read_in;
  /* control.vhdl:162:70  */
  assign n27276_o = n27272_o & n27275_o;
  assign n27278_o = {gpr_b_read_valid_in, 2'b00};
  /* control.vhdl:162:13  */
  assign n27280_o = n27276_o ? n27278_o : 3'b000;
  /* control.vhdl:162:24  */
  assign n27282_o = tag_regs[29:20];
  /* control.vhdl:162:28  */
  assign n27283_o = n27282_o[0];
  /* control.vhdl:162:53  */
  assign n27284_o = tag_regs[29:20];
  /* control.vhdl:162:57  */
  assign n27285_o = n27284_o[8];
  /* control.vhdl:162:41  */
  assign n27286_o = n27283_o & n27285_o;
  /* control.vhdl:162:82  */
  assign n27287_o = tag_regs[29:20];
  /* control.vhdl:162:86  */
  assign n27288_o = n27287_o[7:1];
  /* control.vhdl:162:90  */
  assign n27289_o = n27288_o == gpr_b_read_in;
  /* control.vhdl:162:70  */
  assign n27290_o = n27286_o & n27289_o;
  assign n27292_o = {gpr_b_read_valid_in, 2'b01};
  /* control.vhdl:162:13  */
  assign n27293_o = n27290_o ? n27292_o : n27280_o;
  /* control.vhdl:162:24  */
  assign n27294_o = tag_regs[19:10];
  /* control.vhdl:162:28  */
  assign n27295_o = n27294_o[0];
  /* control.vhdl:162:53  */
  assign n27296_o = tag_regs[19:10];
  /* control.vhdl:162:57  */
  assign n27297_o = n27296_o[8];
  /* control.vhdl:162:41  */
  assign n27298_o = n27295_o & n27297_o;
  /* control.vhdl:162:82  */
  assign n27299_o = tag_regs[19:10];
  /* control.vhdl:162:86  */
  assign n27300_o = n27299_o[7:1];
  /* control.vhdl:162:90  */
  assign n27301_o = n27300_o == gpr_b_read_in;
  /* control.vhdl:162:70  */
  assign n27302_o = n27298_o & n27301_o;
  assign n27304_o = {gpr_b_read_valid_in, 2'b10};
  /* control.vhdl:162:13  */
  assign n27305_o = n27302_o ? n27304_o : n27293_o;
  /* control.vhdl:162:24  */
  assign n27306_o = tag_regs[9:0];
  /* control.vhdl:162:28  */
  assign n27307_o = n27306_o[0];
  /* control.vhdl:162:53  */
  assign n27308_o = tag_regs[9:0];
  /* control.vhdl:162:57  */
  assign n27309_o = n27308_o[8];
  /* control.vhdl:162:41  */
  assign n27310_o = n27307_o & n27309_o;
  /* control.vhdl:162:82  */
  assign n27311_o = tag_regs[9:0];
  /* control.vhdl:162:86  */
  assign n27312_o = n27311_o[7:1];
  /* control.vhdl:162:90  */
  assign n27313_o = n27312_o == gpr_b_read_in;
  /* control.vhdl:162:70  */
  assign n27314_o = n27310_o & n27313_o;
  assign n27316_o = {gpr_b_read_valid_in, 2'b11};
  /* control.vhdl:162:13  */
  assign n27317_o = n27314_o ? n27316_o : n27305_o;
  /* common.vhdl:785:21  */
  assign n27323_o = n27317_o[2];
  /* common.vhdl:785:42  */
  assign n27324_o = n26964_o[2];
  /* common.vhdl:785:33  */
  assign n27325_o = n27323_o & n27324_o;
  /* common.vhdl:785:63  */
  assign n27326_o = n27317_o[1:0];
  /* common.vhdl:785:67  */
  assign n27327_o = {30'b0, n27326_o};  //  uext
  /* common.vhdl:785:74  */
  assign n27328_o = n26964_o[1:0];
  /* common.vhdl:785:67  */
  assign n27329_o = {30'b0, n27328_o};  //  uext
  /* common.vhdl:785:67  */
  assign n27330_o = n27327_o == n27329_o;
  /* common.vhdl:785:54  */
  assign n27331_o = n27325_o & n27330_o;
  assign n27333_o = n27316_o[2];
  assign n27334_o = n27304_o[2];
  assign n27335_o = n27292_o[2];
  assign n27336_o = n27278_o[2];
  assign n27337_o = n27279_o[2];
  /* control.vhdl:162:13  */
  assign n27338_o = n27276_o ? n27336_o : n27337_o;
  /* control.vhdl:162:13  */
  assign n27339_o = n27290_o ? n27335_o : n27338_o;
  /* control.vhdl:162:13  */
  assign n27340_o = n27302_o ? n27334_o : n27339_o;
  /* control.vhdl:162:13  */
  assign n27341_o = n27314_o ? n27333_o : n27340_o;
  /* control.vhdl:167:9  */
  assign n27342_o = n27331_o ? 1'b0 : n27341_o;
  assign n27343_o = n27316_o[1:0];
  assign n27344_o = n27304_o[1:0];
  assign n27345_o = n27292_o[1:0];
  assign n27346_o = n27278_o[1:0];
  assign n27347_o = n27279_o[1:0];
  /* control.vhdl:162:13  */
  assign n27348_o = n27276_o ? n27346_o : n27347_o;
  /* control.vhdl:162:13  */
  assign n27349_o = n27290_o ? n27345_o : n27348_o;
  /* control.vhdl:162:13  */
  assign n27350_o = n27302_o ? n27344_o : n27349_o;
  /* control.vhdl:162:13  */
  assign n27351_o = n27314_o ? n27343_o : n27350_o;
  /* control.vhdl:172:24  */
  assign n27352_o = tag_regs[39:30];
  /* control.vhdl:172:28  */
  assign n27353_o = n27352_o[0];
  /* control.vhdl:172:53  */
  assign n27354_o = tag_regs[39:30];
  /* control.vhdl:172:57  */
  assign n27355_o = n27354_o[8];
  /* control.vhdl:172:41  */
  assign n27356_o = n27353_o & n27355_o;
  /* control.vhdl:172:82  */
  assign n27357_o = tag_regs[39:30];
  /* control.vhdl:172:86  */
  assign n27358_o = n27357_o[7:1];
  /* control.vhdl:172:90  */
  assign n27359_o = n27358_o == gpr_c_read_in;
  /* control.vhdl:172:70  */
  assign n27360_o = n27356_o & n27359_o;
  assign n27362_o = {gpr_c_read_valid_in, 2'b00};
  /* control.vhdl:172:13  */
  assign n27364_o = n27360_o ? n27362_o : 3'b000;
  /* control.vhdl:172:24  */
  assign n27366_o = tag_regs[29:20];
  /* control.vhdl:172:28  */
  assign n27367_o = n27366_o[0];
  /* control.vhdl:172:53  */
  assign n27368_o = tag_regs[29:20];
  /* control.vhdl:172:57  */
  assign n27369_o = n27368_o[8];
  /* control.vhdl:172:41  */
  assign n27370_o = n27367_o & n27369_o;
  /* control.vhdl:172:82  */
  assign n27371_o = tag_regs[29:20];
  /* control.vhdl:172:86  */
  assign n27372_o = n27371_o[7:1];
  /* control.vhdl:172:90  */
  assign n27373_o = n27372_o == gpr_c_read_in;
  /* control.vhdl:172:70  */
  assign n27374_o = n27370_o & n27373_o;
  assign n27376_o = {gpr_c_read_valid_in, 2'b01};
  /* control.vhdl:172:13  */
  assign n27377_o = n27374_o ? n27376_o : n27364_o;
  /* control.vhdl:172:24  */
  assign n27378_o = tag_regs[19:10];
  /* control.vhdl:172:28  */
  assign n27379_o = n27378_o[0];
  /* control.vhdl:172:53  */
  assign n27380_o = tag_regs[19:10];
  /* control.vhdl:172:57  */
  assign n27381_o = n27380_o[8];
  /* control.vhdl:172:41  */
  assign n27382_o = n27379_o & n27381_o;
  /* control.vhdl:172:82  */
  assign n27383_o = tag_regs[19:10];
  /* control.vhdl:172:86  */
  assign n27384_o = n27383_o[7:1];
  /* control.vhdl:172:90  */
  assign n27385_o = n27384_o == gpr_c_read_in;
  /* control.vhdl:172:70  */
  assign n27386_o = n27382_o & n27385_o;
  assign n27388_o = {gpr_c_read_valid_in, 2'b10};
  /* control.vhdl:172:13  */
  assign n27389_o = n27386_o ? n27388_o : n27377_o;
  /* control.vhdl:172:24  */
  assign n27390_o = tag_regs[9:0];
  /* control.vhdl:172:28  */
  assign n27391_o = n27390_o[0];
  /* control.vhdl:172:53  */
  assign n27392_o = tag_regs[9:0];
  /* control.vhdl:172:57  */
  assign n27393_o = n27392_o[8];
  /* control.vhdl:172:41  */
  assign n27394_o = n27391_o & n27393_o;
  /* control.vhdl:172:82  */
  assign n27395_o = tag_regs[9:0];
  /* control.vhdl:172:86  */
  assign n27396_o = n27395_o[7:1];
  /* control.vhdl:172:90  */
  assign n27397_o = n27396_o == gpr_c_read_in;
  /* control.vhdl:172:70  */
  assign n27398_o = n27394_o & n27397_o;
  assign n27400_o = {gpr_c_read_valid_in, 2'b11};
  /* control.vhdl:172:13  */
  assign n27401_o = n27398_o ? n27400_o : n27389_o;
  /* common.vhdl:785:21  */
  assign n27407_o = n27401_o[2];
  /* common.vhdl:785:42  */
  assign n27408_o = n26964_o[2];
  /* common.vhdl:785:33  */
  assign n27409_o = n27407_o & n27408_o;
  /* common.vhdl:785:63  */
  assign n27410_o = n27401_o[1:0];
  /* common.vhdl:785:67  */
  assign n27411_o = {30'b0, n27410_o};  //  uext
  /* common.vhdl:785:74  */
  assign n27412_o = n26964_o[1:0];
  /* common.vhdl:785:67  */
  assign n27413_o = {30'b0, n27412_o};  //  uext
  /* common.vhdl:785:67  */
  assign n27414_o = n27411_o == n27413_o;
  /* common.vhdl:785:54  */
  assign n27415_o = n27409_o & n27414_o;
  assign n27417_o = n27400_o[2];
  assign n27418_o = n27388_o[2];
  assign n27419_o = n27376_o[2];
  assign n27420_o = n27362_o[2];
  assign n27421_o = n27363_o[2];
  /* control.vhdl:172:13  */
  assign n27422_o = n27360_o ? n27420_o : n27421_o;
  /* control.vhdl:172:13  */
  assign n27423_o = n27374_o ? n27419_o : n27422_o;
  /* control.vhdl:172:13  */
  assign n27424_o = n27386_o ? n27418_o : n27423_o;
  /* control.vhdl:172:13  */
  assign n27425_o = n27398_o ? n27417_o : n27424_o;
  /* control.vhdl:177:9  */
  assign n27426_o = n27415_o ? 1'b0 : n27425_o;
  assign n27427_o = n27400_o[1:0];
  assign n27428_o = n27388_o[1:0];
  assign n27429_o = n27376_o[1:0];
  assign n27430_o = n27362_o[1:0];
  assign n27431_o = n27363_o[1:0];
  /* control.vhdl:172:13  */
  assign n27432_o = n27360_o ? n27430_o : n27431_o;
  /* control.vhdl:172:13  */
  assign n27433_o = n27374_o ? n27429_o : n27432_o;
  /* control.vhdl:172:13  */
  assign n27434_o = n27386_o ? n27428_o : n27433_o;
  /* control.vhdl:172:13  */
  assign n27435_o = n27398_o ? n27427_o : n27434_o;
  /* common.vhdl:785:21  */
  assign n27441_o = n26965_o[2];
  assign n27442_o = {n27258_o, n27267_o};
  /* common.vhdl:785:42  */
  assign n27443_o = n27442_o[2];
  /* common.vhdl:785:33  */
  assign n27444_o = n27441_o & n27443_o;
  /* common.vhdl:785:63  */
  assign n27445_o = n26965_o[1:0];
  /* common.vhdl:785:67  */
  assign n27446_o = {30'b0, n27445_o};  //  uext
  assign n27447_o = {n27258_o, n27267_o};
  /* common.vhdl:785:74  */
  assign n27448_o = n27447_o[1:0];
  /* common.vhdl:785:67  */
  assign n27449_o = {30'b0, n27448_o};  //  uext
  /* common.vhdl:785:67  */
  assign n27450_o = n27446_o == n27449_o;
  /* common.vhdl:785:54  */
  assign n27451_o = n27444_o & n27450_o;
  /* control.vhdl:182:23  */
  assign n27453_o = 1'b1 & n27451_o;
  /* control.vhdl:182:9  */
  assign n27456_o = n27453_o ? 1'b1 : 1'b0;
  /* common.vhdl:785:21  */
  assign n27463_o = n26965_o[2];
  assign n27464_o = {n27342_o, n27351_o};
  /* common.vhdl:785:42  */
  assign n27465_o = n27464_o[2];
  /* common.vhdl:785:33  */
  assign n27466_o = n27463_o & n27465_o;
  /* common.vhdl:785:63  */
  assign n27467_o = n26965_o[1:0];
  /* common.vhdl:785:67  */
  assign n27468_o = {30'b0, n27467_o};  //  uext
  assign n27469_o = {n27342_o, n27351_o};
  /* common.vhdl:785:74  */
  assign n27470_o = n27469_o[1:0];
  /* common.vhdl:785:67  */
  assign n27471_o = {30'b0, n27470_o};  //  uext
  /* common.vhdl:785:67  */
  assign n27472_o = n27468_o == n27471_o;
  /* common.vhdl:785:54  */
  assign n27473_o = n27466_o & n27472_o;
  /* control.vhdl:186:23  */
  assign n27475_o = 1'b1 & n27473_o;
  /* control.vhdl:186:9  */
  assign n27478_o = n27475_o ? 1'b1 : 1'b0;
  /* common.vhdl:785:21  */
  assign n27485_o = n26965_o[2];
  assign n27486_o = {n27426_o, n27435_o};
  /* common.vhdl:785:42  */
  assign n27487_o = n27486_o[2];
  /* common.vhdl:785:33  */
  assign n27488_o = n27485_o & n27487_o;
  /* common.vhdl:785:63  */
  assign n27489_o = n26965_o[1:0];
  /* common.vhdl:785:67  */
  assign n27490_o = {30'b0, n27489_o};  //  uext
  assign n27491_o = {n27426_o, n27435_o};
  /* common.vhdl:785:74  */
  assign n27492_o = n27491_o[1:0];
  /* common.vhdl:785:67  */
  assign n27493_o = {30'b0, n27492_o};  //  uext
  /* common.vhdl:785:67  */
  assign n27494_o = n27490_o == n27493_o;
  /* common.vhdl:785:54  */
  assign n27495_o = n27488_o & n27494_o;
  /* control.vhdl:190:23  */
  assign n27497_o = 1'b1 & n27495_o;
  /* control.vhdl:190:9  */
  assign n27500_o = n27497_o ? 1'b1 : 1'b0;
  assign n27502_o = {n27258_o, n27267_o};
  /* control.vhdl:198:33  */
  assign n27503_o = n27502_o[2];
  /* control.vhdl:198:43  */
  assign n27504_o = ~n27456_o;
  /* control.vhdl:198:39  */
  assign n27505_o = n27503_o & n27504_o;
  assign n27506_o = {n27342_o, n27351_o};
  /* control.vhdl:199:33  */
  assign n27507_o = n27506_o[2];
  /* control.vhdl:199:43  */
  assign n27508_o = ~n27478_o;
  /* control.vhdl:199:39  */
  assign n27509_o = n27507_o & n27508_o;
  /* control.vhdl:198:54  */
  assign n27510_o = n27505_o | n27509_o;
  assign n27511_o = {n27426_o, n27435_o};
  /* control.vhdl:200:33  */
  assign n27512_o = n27511_o[2];
  /* control.vhdl:200:43  */
  assign n27513_o = ~n27500_o;
  /* control.vhdl:200:39  */
  assign n27514_o = n27512_o & n27513_o;
  /* control.vhdl:199:54  */
  assign n27515_o = n27510_o | n27514_o;
  /* control.vhdl:204:42  */
  assign n27516_o = ~deferred;
  /* control.vhdl:204:38  */
  assign n27517_o = n27702_o & n27516_o;
  /* control.vhdl:205:22  */
  assign n27518_o = instr_tag[2];
  /* control.vhdl:206:35  */
  assign n27519_o = {30'b0, curr_tag};  //  uext
  /* control.vhdl:206:35  */
  assign n27521_o = n27519_o + 32'b00000000000000000000000000000001;
  assign n27522_o = n27521_o[1:0];
  /* control.vhdl:205:9  */
  assign n27524_o = n27518_o ? n27522_o : curr_tag;
  /* control.vhdl:213:49  */
  assign n27526_o = 2'b11 - curr_cr_tag;
  /* control.vhdl:213:62  */
  assign n27529_o = n27729_o[9];
  /* control.vhdl:213:36  */
  assign n27530_o = cr_read_in & n27529_o;
  assign n27536_o = {n27530_o, curr_cr_tag};
  /* common.vhdl:785:21  */
  assign n27537_o = n27536_o[2];
  /* common.vhdl:785:42  */
  assign n27538_o = n26964_o[2];
  /* common.vhdl:785:33  */
  assign n27539_o = n27537_o & n27538_o;
  assign n27540_o = {n27530_o, curr_cr_tag};
  /* common.vhdl:785:63  */
  assign n27541_o = n27540_o[1:0];
  /* common.vhdl:785:67  */
  assign n27542_o = {30'b0, n27541_o};  //  uext
  /* common.vhdl:785:74  */
  assign n27543_o = n26964_o[1:0];
  /* common.vhdl:785:67  */
  assign n27544_o = {30'b0, n27543_o};  //  uext
  /* common.vhdl:785:67  */
  assign n27545_o = n27542_o == n27544_o;
  /* common.vhdl:785:54  */
  assign n27546_o = n27539_o & n27545_o;
  /* control.vhdl:214:9  */
  assign n27548_o = n27546_o ? 1'b0 : n27530_o;
  /* common.vhdl:785:21  */
  assign n27554_o = n26966_o[2];
  assign n27555_o = {n27548_o, curr_cr_tag};
  /* common.vhdl:785:42  */
  assign n27556_o = n27555_o[2];
  /* common.vhdl:785:33  */
  assign n27557_o = n27554_o & n27556_o;
  /* common.vhdl:785:63  */
  assign n27558_o = n26966_o[1:0];
  /* common.vhdl:785:67  */
  assign n27559_o = {30'b0, n27558_o};  //  uext
  assign n27560_o = {n27548_o, curr_cr_tag};
  /* common.vhdl:785:74  */
  assign n27561_o = n27560_o[1:0];
  /* common.vhdl:785:67  */
  assign n27562_o = {30'b0, n27561_o};  //  uext
  /* common.vhdl:785:67  */
  assign n27563_o = n27559_o == n27562_o;
  /* common.vhdl:785:54  */
  assign n27564_o = n27557_o & n27563_o;
  /* control.vhdl:218:23  */
  assign n27566_o = 1'b1 & n27564_o;
  /* control.vhdl:218:9  */
  assign n27569_o = n27566_o ? 1'b1 : 1'b0;
  assign n27571_o = {n27548_o, curr_cr_tag};
  /* control.vhdl:223:32  */
  assign n27572_o = n27571_o[2];
  /* control.vhdl:223:42  */
  assign n27573_o = ~n27569_o;
  /* control.vhdl:223:38  */
  assign n27574_o = n27572_o & n27573_o;
  /* control.vhdl:234:35  */
  assign n27589_o = ~flush_in;
  /* control.vhdl:234:31  */
  assign n27590_o = valid_in & n27589_o;
  /* control.vhdl:239:27  */
  assign n27592_o = n26964_o[2];
  /* control.vhdl:240:40  */
  assign n27593_o = r_int[5:2];
  /* control.vhdl:240:52  */
  assign n27594_o = {{28{n27593_o[3]}}, n27593_o}; // sext
  /* control.vhdl:240:52  */
  assign n27596_o = n27594_o - 32'b00000000000000000000000000000001;
  /* control.vhdl:240:13  */
  assign n27597_o = n27596_o[3:0];  // trunc
  assign n27598_o = r_int[5:2];
  /* control.vhdl:239:9  */
  assign n27599_o = n27592_o ? n27597_o : n27598_o;
  /* control.vhdl:237:9  */
  assign n27600_o = flush_in ? 4'b0000 : n27599_o;
  assign n27601_o = r_int[1:0];
  /* control.vhdl:242:18  */
  assign n27602_o = r_int[5:2];
  /* control.vhdl:242:30  */
  assign n27603_o = {{28{n27602_o[3]}}, n27602_o}; // sext
  /* control.vhdl:242:30  */
  assign n27605_o = $signed(n27603_o) >= $signed(32'b00000000000000000000000000000100);
  /* control.vhdl:242:9  */
  assign n27607_o = n27605_o ? 1'b0 : n27590_o;
  /* control.vhdl:242:9  */
  assign n27610_o = n27605_o ? 1'b1 : 1'b0;
  assign n27613_o = {n27600_o, n27601_o};
  /* control.vhdl:247:9  */
  assign n27614_o = rst ? 6'b000000 : n27613_o;
  /* control.vhdl:247:9  */
  assign n27616_o = rst ? 1'b0 : n27607_o;
  /* control.vhdl:254:41  */
  assign n27617_o = n27614_o[5:2];
  /* control.vhdl:254:53  */
  assign n27618_o = {{28{n27617_o[3]}}, n27617_o}; // sext
  /* control.vhdl:254:53  */
  assign n27620_o = n27618_o == 32'b00000000000000000000000000000000;
  /* control.vhdl:254:31  */
  assign n27621_o = stop_mark_in & n27620_o;
  /* control.vhdl:254:9  */
  assign n27624_o = n27621_o ? 1'b1 : 1'b0;
  /* control.vhdl:260:20  */
  assign n27626_o = r_int[1:0];
  /* control.vhdl:264:34  */
  assign n27627_o = n27614_o[5:2];
  /* control.vhdl:264:46  */
  assign n27628_o = {{28{n27627_o[3]}}, n27627_o}; // sext
  /* control.vhdl:264:46  */
  assign n27630_o = n27628_o != 32'b00000000000000000000000000000000;
  /* control.vhdl:264:25  */
  assign n27633_o = n27630_o ? 2'b01 : 2'b10;
  /* control.vhdl:264:25  */
  assign n27635_o = n27630_o ? 1'b1 : n27610_o;
  /* control.vhdl:273:52  */
  assign n27636_o = gpr_tag_stall | cr_tag_stall;
  assign n27637_o = n27612_o[1:0];
  assign n27638_o = n27613_o[1:0];
  /* control.vhdl:247:9  */
  assign n27639_o = rst ? n27637_o : n27638_o;
  /* control.vhdl:263:21  */
  assign n27640_o = sgl_pipe_in ? n27633_o : n27639_o;
  /* control.vhdl:263:21  */
  assign n27641_o = sgl_pipe_in ? n27635_o : n27636_o;
  assign n27642_o = n27612_o[1:0];
  assign n27643_o = n27613_o[1:0];
  /* control.vhdl:247:9  */
  assign n27644_o = rst ? n27642_o : n27643_o;
  /* control.vhdl:262:17  */
  assign n27645_o = n27616_o ? n27640_o : n27644_o;
  /* control.vhdl:262:17  */
  assign n27646_o = n27616_o ? n27641_o : n27610_o;
  /* control.vhdl:261:13  */
  assign n27648_o = n27626_o == 2'b00;
  /* control.vhdl:278:26  */
  assign n27649_o = n27614_o[5:2];
  /* control.vhdl:278:38  */
  assign n27650_o = {{28{n27649_o[3]}}, n27649_o}; // sext
  /* control.vhdl:278:38  */
  assign n27652_o = n27650_o == 32'b00000000000000000000000000000000;
  assign n27654_o = n27612_o[1:0];
  assign n27655_o = n27613_o[1:0];
  /* control.vhdl:247:9  */
  assign n27656_o = rst ? n27654_o : n27655_o;
  /* control.vhdl:278:17  */
  assign n27657_o = n27652_o ? 2'b10 : n27656_o;
  /* control.vhdl:278:17  */
  assign n27659_o = n27652_o ? n27610_o : 1'b1;
  /* control.vhdl:277:13  */
  assign n27661_o = n27626_o == 2'b01;
  /* control.vhdl:286:26  */
  assign n27662_o = n27614_o[5:2];
  /* control.vhdl:286:38  */
  assign n27663_o = {{28{n27662_o[3]}}, n27662_o}; // sext
  /* control.vhdl:286:38  */
  assign n27665_o = n27663_o == 32'b00000000000000000000000000000000;
  assign n27667_o = n27612_o[5:2];
  assign n27668_o = n27613_o[5:2];
  /* control.vhdl:247:9  */
  assign n27669_o = rst ? n27667_o : n27668_o;
  assign n27670_o = {n27669_o, 2'b00};
  /* control.vhdl:291:38  */
  assign n27671_o = n27670_o[5:2];
  /* control.vhdl:291:50  */
  assign n27672_o = {{28{n27671_o[3]}}, n27671_o}; // sext
  /* control.vhdl:291:50  */
  assign n27674_o = n27672_o != 32'b00000000000000000000000000000000;
  /* control.vhdl:291:29  */
  assign n27677_o = n27674_o ? 2'b01 : 2'b10;
  /* control.vhdl:291:29  */
  assign n27679_o = n27674_o ? 1'b1 : n27610_o;
  /* control.vhdl:300:56  */
  assign n27680_o = gpr_tag_stall | cr_tag_stall;
  /* control.vhdl:289:21  */
  assign n27681_o = n27683_o ? n27677_o : 2'b00;
  /* control.vhdl:290:25  */
  assign n27682_o = sgl_pipe_in ? n27679_o : n27680_o;
  /* control.vhdl:289:21  */
  assign n27683_o = n27616_o & sgl_pipe_in;
  /* control.vhdl:289:21  */
  assign n27684_o = n27616_o ? n27682_o : n27610_o;
  assign n27685_o = n27612_o[1:0];
  assign n27686_o = n27613_o[1:0];
  /* control.vhdl:247:9  */
  assign n27687_o = rst ? n27685_o : n27686_o;
  /* control.vhdl:286:17  */
  assign n27688_o = n27665_o ? n27681_o : n27687_o;
  /* control.vhdl:286:17  */
  assign n27690_o = n27665_o ? n27684_o : 1'b1;
  /* control.vhdl:285:13  */
  assign n27692_o = n27626_o == 2'b10;
  assign n27693_o = {n27692_o, n27661_o, n27648_o};
  /* control.vhdl:260:9  */
  always @*
    case (n27693_o)
      3'b100: n27695_o = n27688_o;
      3'b010: n27695_o = n27657_o;
      3'b001: n27695_o = n27645_o;
      default: n27695_o = 2'bX;
    endcase
  assign n27696_o = n27612_o[5:2];
  assign n27697_o = n27613_o[5:2];
  /* control.vhdl:247:9  */
  assign n27698_o = rst ? n27696_o : n27697_o;
  /* control.vhdl:260:9  */
  always @*
    case (n27693_o)
      3'b100: n27700_o = n27690_o;
      3'b010: n27700_o = n27659_o;
      3'b001: n27700_o = n27646_o;
      default: n27700_o = 1'bX;
    endcase
  /* control.vhdl:308:9  */
  assign n27702_o = n27700_o ? 1'b0 : n27616_o;
  /* control.vhdl:312:47  */
  assign n27703_o = gpr_write_valid_in & n27702_o;
  /* control.vhdl:313:39  */
  assign n27704_o = cr_write_in & n27702_o;
  /* control.vhdl:315:41  */
  assign n27705_o = ~deferred;
  /* control.vhdl:315:28  */
  assign n27706_o = n27702_o & n27705_o;
  assign n27707_o = {n27698_o, n27695_o};
  /* control.vhdl:316:40  */
  assign n27708_o = n27707_o[5:2];
  /* control.vhdl:316:52  */
  assign n27709_o = {{28{n27708_o[3]}}, n27708_o}; // sext
  /* control.vhdl:316:52  */
  assign n27711_o = n27709_o + 32'b00000000000000000000000000000001;
  /* control.vhdl:316:13  */
  assign n27712_o = n27711_o[3:0];  // trunc
  /* control.vhdl:315:9  */
  assign n27713_o = n27706_o ? n27712_o : n27698_o;
  /* control.vhdl:321:32  */
  assign n27714_o = n27700_o | deferred;
  assign n27715_o = {n27713_o, n27695_o};
  /* control.vhdl:93:9  */
  always @(posedge clk)
    n27719_q <= rin_int;
  initial
    n27719_q = 6'b000000;
  /* control.vhdl:93:9  */
  always @(posedge clk)
    n27720_q <= n27166_o;
  /* control.vhdl:93:9  */
  assign n27721_o = {n27517_o, curr_tag};
  /* control.vhdl:93:9  */
  always @(posedge clk)
    n27722_q <= n27162_o;
  /* control.vhdl:93:9  */
  always @(posedge clk)
    n27723_q <= n27164_o;
  assign n27724_o = tag_regs[9:0];
  assign n27725_o = tag_regs[19:10];
  assign n27726_o = tag_regs[29:20];
  assign n27727_o = tag_regs[39:30];
  /* control.vhdl:213:48  */
  assign n27728_o = n27526_o[1:0];
  /* control.vhdl:213:48  */
  always @*
    case (n27728_o)
      2'b00: n27729_o = n27724_o;
      2'b01: n27729_o = n27725_o;
      2'b10: n27729_o = n27726_o;
      2'b11: n27729_o = n27727_o;
    endcase
endmodule

module cache_ram_5_64_1489f923c4dca729178b3e3233458550d8dddf29
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  clk,
   input  rd_en,
   input  [4:0] rd_addr,
   input  [7:0] wr_sel,
   input  [4:0] wr_addr,
   input  [63:0] wr_data,
   output [63:0] rd_data);
  wire wr_enable;
  wire [63:0] rd_data0_tmp;
  wire [63:0] rd_data0_saved;
  wire [63:0] rd_data0;
  wire rd_en_prev;
  wire n26951_o;
  wire [63:0] cache_ram_0_Do0;
  wire [63:0] cache_ram_0_Do1;
  wire [63:0] n26960_o;
  wire [63:0] n26961_o;
  reg [63:0] n26962_q;
  reg n26963_q;
  assign rd_data = rd_data0;
  /* asic/cache_ram.vhdl:44:12  */
  assign wr_enable = n26951_o; // (signal)
  /* asic/cache_ram.vhdl:45:12  */
  assign rd_data0_tmp = cache_ram_0_Do1; // (signal)
  /* asic/cache_ram.vhdl:46:12  */
  assign rd_data0_saved = n26962_q; // (signal)
  /* asic/cache_ram.vhdl:47:12  */
  assign rd_data0 = n26960_o; // (signal)
  /* asic/cache_ram.vhdl:48:12  */
  assign rd_en_prev = n26963_q; // (signal)
  /* asic/cache_ram.vhdl:54:18  */
  assign n26951_o = |(wr_sel);
  /* asic/cache_ram.vhdl:56:5  */
  RAM32_1RW1R cache_ram_0 (
`ifdef USE_POWER_PINS
    .VPWR(vccd1),
    .VGND(vssd1),
`endif
    .CLK(clk),
    .EN0(wr_enable),
    .A0(wr_addr),
    .WE0(wr_sel),
    .Di0(wr_data),
    .EN1(rd_en),
    .A1(rd_addr),
    .Do0(),
    .Do1(cache_ram_0_Do1));
  /* asic/cache_ram.vhdl:82:30  */
  assign n26960_o = rd_en_prev ? rd_data0_tmp : rd_data0_saved;
  /* asic/cache_ram.vhdl:75:9  */
  assign n26961_o = rd_en_prev ? rd_data0_tmp : rd_data0_saved;
  /* asic/cache_ram.vhdl:75:9  */
  always @(posedge clk)
    n26962_q <= n26961_o;
  /* asic/cache_ram.vhdl:75:9  */
  always @(posedge clk)
    n26963_q <= rd_en;
endmodule

module main_bram_64_9_4096_a75adb9e07879fb6c63b494abe06e3f9a6bb2ed9
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  clk,
   input  [8:0] addr,
   input  [63:0] din,
   input  [7:0] sel,
   input  re,
   input  we,
   output [63:0] dout);
  wire [7:0] sel_qual;
  wire [63:0] obuf;
  wire [7:0] n26941_o;
  wire [63:0] memory_0_Do0;
  wire n26943_o;
  reg [63:0] n26949_q;
  assign dout = n26949_q;
  /* asic/main_bram.vhdl:49:29  */
  assign sel_qual = n26941_o; // (signal)
  /* asic/main_bram.vhdl:37:12  */
  assign obuf = memory_0_Do0; // (signal)
  /* asic/main_bram.vhdl:44:21  */
  assign n26941_o = we ? sel : 8'b00000000;
  /* asic/main_bram.vhdl:46:5  */
  RAM512 memory_0 (
`ifdef USE_POWER_PINS
    .VPWR(vccd1),
    .VGND(vssd1),
`endif
    .CLK(clk),
    .WE0(sel_qual),
    .EN0(n26943_o),
    .Di0(din),
    .A0(addr),
    .Do0(memory_0_Do0));
  /* asic/main_bram.vhdl:50:24  */
  assign n26943_o = re | we;
  /* asic/main_bram.vhdl:59:9  */
  always @(posedge clk)
    n26949_q <= obuf;
endmodule

module spi_rxtx_4_1
  (input  clk,
   input  rst,
   input  [7:0] clk_div_i,
   input  cmd_valid_i,
   input  [2:0] cmd_mode_i,
   input  [2:0] cmd_clks_i,
   input  [7:0] cmd_txd_i,
   input  [3:0] sdat_i,
   output cmd_ready_o,
   output [7:0] d_rxd_o,
   output d_ack_o,
   output bus_idle_o,
   output sck,
   output [3:0] sdat_o,
   output [3:0] sdat_oe);
  wire sck_0;
  wire sck_1;
  wire [7:0] clk_div;
  wire sck_send;
  wire sck_recv;
  wire [2:0] cmd_mode;
  wire [7:0] oreg;
  wire [3:0] dat_i_l;
  wire dat_ack_l;
  reg sck_recv_d;
  reg [7:0] ireg;
  wire [2:0] bit_count;
  wire next_cmd;
  wire start_cmd;
  wire end_cmd;
  reg state;
  reg [7:0] sck_gen_counter;
  wire [31:0] n26629_o;
  wire [31:0] n26630_o;
  wire n26631_o;
  wire n26632_o;
  wire n26633_o;
  wire [31:0] n26634_o;
  wire [31:0] n26636_o;
  wire [7:0] n26637_o;
  wire n26638_o;
  wire [7:0] n26639_o;
  wire n26641_o;
  wire n26643_o;
  wire [7:0] n26645_o;
  wire n26647_o;
  wire [7:0] n26651_o;
  wire n26653_o;
  wire n26655_o;
  wire [7:0] n26657_o;
  wire n26659_o;
  wire n26660_o;
  wire n26661_o;
  wire n26662_o;
  wire n26663_o;
  wire n26665_o;
  reg [7:0] n26673_q;
  wire n26676_o;
  wire n26677_o;
  wire n26678_o;
  wire n26680_o;
  wire n26681_o;
  wire n26682_o;
  wire n26685_o;
  wire n26686_o;
  wire n26691_o;
  wire [2:0] n26692_o;
  wire n26694_o;
  wire [2:0] n26696_o;
  wire n26698_o;
  wire n26705_o;
  wire [2:0] n26707_o;
  wire [2:0] n26708_o;
  wire [2:0] n26710_o;
  wire [2:0] n26711_o;
  wire [2:0] n26713_o;
  wire n26723_o;
  wire n26724_o;
  wire [6:0] n26725_o;
  wire [7:0] n26727_o;
  wire [1:0] n26733_o;
  wire n26735_o;
  wire [5:0] n26736_o;
  wire [7:0] n26738_o;
  wire [3:0] n26739_o;
  wire [7:0] n26741_o;
  wire [7:0] n26742_o;
  wire [7:0] n26743_o;
  wire [7:0] n26744_o;
  wire [7:0] n26745_o;
  wire n26748_o;
  wire n26749_o;
  wire n26750_o;
  wire n26751_o;
  wire n26755_o;
  wire [1:0] n26761_o;
  wire n26763_o;
  wire n26765_o;
  wire n26771_o;
  wire n26772_o;
  wire n26774_o;
  wire n26775_o;
  wire n26778_o;
  wire [1:0] n26784_o;
  wire n26786_o;
  wire n26788_o;
  wire n26794_o;
  wire n26795_o;
  wire n26797_o;
  wire n26798_o;
  wire n26801_o;
  wire [1:0] n26807_o;
  wire n26809_o;
  wire n26811_o;
  wire n26817_o;
  wire n26818_o;
  wire n26820_o;
  wire [1:0] n26826_o;
  wire n26828_o;
  wire n26830_o;
  wire n26836_o;
  wire n26837_o;
  wire n26839_o;
  wire n26840_o;
  wire n26843_o;
  wire n26849_o;
  wire n26850_o;
  wire n26856_o;
  wire n26857_o;
  wire n26859_o;
  wire n26861_o;
  wire n26862_o;
  wire n26872_o;
  wire n26874_o;
  wire n26876_o;
  wire n26877_o;
  wire n26878_o;
  wire n26879_o;
  wire n26881_o;
  wire [1:0] n26887_o;
  wire n26889_o;
  wire [5:0] n26890_o;
  wire n26891_o;
  wire [6:0] n26892_o;
  wire n26893_o;
  wire [7:0] n26894_o;
  wire [1:0] n26900_o;
  wire n26902_o;
  wire [3:0] n26903_o;
  wire n26904_o;
  wire [4:0] n26905_o;
  wire n26906_o;
  wire [5:0] n26907_o;
  wire n26908_o;
  wire [6:0] n26909_o;
  wire n26910_o;
  wire [7:0] n26911_o;
  wire [6:0] n26912_o;
  wire n26913_o;
  wire [7:0] n26914_o;
  wire [7:0] n26915_o;
  wire [7:0] n26916_o;
  reg n26923_q;
  reg n26924_q;
  reg [7:0] n26925_q;
  reg n26926_q;
  reg n26927_q;
  reg [2:0] n26928_q;
  reg [7:0] n26929_q;
  reg [3:0] n26930_q;
  reg n26931_q;
  reg n26932_q;
  wire [7:0] n26933_o;
  reg [7:0] n26934_q;
  reg [2:0] n26935_q;
  reg n26936_q;
  reg n26937_q;
  wire [3:0] n26938_o;
  wire [3:0] n26939_o;
  assign cmd_ready_o = next_cmd;
  assign d_rxd_o = ireg;
  assign d_ack_o = n26937_q;
  assign bus_idle_o = n26686_o;
  assign sck = sck_1;
  assign sdat_o = n26938_o;
  assign sdat_oe = n26939_o;
  /* spi_rxtx.vhdl:98:12  */
  assign sck_0 = n26923_q; // (signal)
  /* spi_rxtx.vhdl:99:12  */
  assign sck_1 = n26924_q; // (signal)
  /* spi_rxtx.vhdl:102:12  */
  assign clk_div = n26925_q; // (signal)
  /* spi_rxtx.vhdl:113:12  */
  assign sck_send = n26926_q; // (signal)
  /* spi_rxtx.vhdl:114:12  */
  assign sck_recv = n26927_q; // (signal)
  /* spi_rxtx.vhdl:117:12  */
  assign cmd_mode = n26928_q; // (signal)
  /* spi_rxtx.vhdl:120:12  */
  assign oreg = n26929_q; // (signal)
  /* spi_rxtx.vhdl:123:12  */
  assign dat_i_l = n26930_q; // (signal)
  /* spi_rxtx.vhdl:126:12  */
  assign dat_ack_l = n26931_q; // (signal)
  /* spi_rxtx.vhdl:129:12  */
  always @*
    sck_recv_d = n26932_q; // (isignal)
  initial
    sck_recv_d = 1'b0;
  /* spi_rxtx.vhdl:132:12  */
  always @*
    ireg = n26934_q; // (isignal)
  initial
    ireg = 8'b00000000;
  /* spi_rxtx.vhdl:135:12  */
  assign bit_count = n26935_q; // (signal)
  /* spi_rxtx.vhdl:138:12  */
  assign next_cmd = n26678_o; // (signal)
  /* spi_rxtx.vhdl:139:12  */
  assign start_cmd = n26680_o; // (signal)
  /* spi_rxtx.vhdl:140:12  */
  assign end_cmd = n26682_o; // (signal)
  /* spi_rxtx.vhdl:160:12  */
  always @*
    state = n26936_q; // (isignal)
  initial
    state = 1'b0;
  /* spi_rxtx.vhdl:171:18  */
  always @*
    sck_gen_counter = n26673_q; // (isignal)
  initial
    sck_gen_counter = 8'b00000000;
  /* spi_rxtx.vhdl:181:27  */
  assign n26629_o = {24'b0, sck_gen_counter};  //  uext
  /* spi_rxtx.vhdl:181:27  */
  assign n26630_o = {24'b0, clk_div};  //  uext
  /* spi_rxtx.vhdl:181:27  */
  assign n26631_o = n26629_o == n26630_o;
  /* spi_rxtx.vhdl:188:26  */
  assign n26632_o = ~sck_0;
  /* spi_rxtx.vhdl:191:29  */
  assign n26633_o = ~sck_0;
  /* spi_rxtx.vhdl:194:36  */
  assign n26634_o = {24'b0, sck_gen_counter};  //  uext
  /* spi_rxtx.vhdl:194:36  */
  assign n26636_o = n26634_o + 32'b00000000000000000000000000000001;
  /* spi_rxtx.vhdl:194:17  */
  assign n26637_o = n26636_o[7:0];  // trunc
  /* spi_rxtx.vhdl:181:13  */
  assign n26638_o = n26631_o ? n26632_o : sck_0;
  /* spi_rxtx.vhdl:181:13  */
  assign n26639_o = n26631_o ? clk_div_i : clk_div;
  /* spi_rxtx.vhdl:181:13  */
  assign n26641_o = n26631_o ? sck_0 : 1'b0;
  /* spi_rxtx.vhdl:181:13  */
  assign n26643_o = n26631_o ? n26633_o : 1'b0;
  /* spi_rxtx.vhdl:181:13  */
  assign n26645_o = n26631_o ? 8'b00000000 : n26637_o;
  /* spi_rxtx.vhdl:174:13  */
  assign n26647_o = rst ? 1'b1 : n26638_o;
  /* spi_rxtx.vhdl:174:13  */
  assign n26651_o = rst ? 8'b00000000 : n26639_o;
  /* spi_rxtx.vhdl:174:13  */
  assign n26653_o = rst ? 1'b0 : n26641_o;
  /* spi_rxtx.vhdl:174:13  */
  assign n26655_o = rst ? 1'b0 : n26643_o;
  /* spi_rxtx.vhdl:174:13  */
  assign n26657_o = rst ? 8'b00000000 : n26645_o;
  /* spi_rxtx.vhdl:203:23  */
  assign n26659_o = state == 1'b1;
  /* spi_rxtx.vhdl:203:42  */
  assign n26660_o = ~end_cmd;
  /* spi_rxtx.vhdl:203:30  */
  assign n26661_o = n26659_o & n26660_o;
  /* spi_rxtx.vhdl:203:68  */
  assign n26662_o = next_cmd & cmd_valid_i;
  /* spi_rxtx.vhdl:203:49  */
  assign n26663_o = n26661_o | n26662_o;
  /* spi_rxtx.vhdl:203:13  */
  assign n26665_o = n26663_o ? sck_0 : 1'b1;
  /* spi_rxtx.vhdl:173:9  */
  always @(posedge clk)
    n26673_q <= n26657_o;
  initial
    n26673_q = 8'b00000000;
  /* spi_rxtx.vhdl:218:56  */
  assign n26676_o = bit_count == 3'b111;
  /* spi_rxtx.vhdl:218:42  */
  assign n26677_o = sck_send & n26676_o;
  /* spi_rxtx.vhdl:218:21  */
  assign n26678_o = n26677_o ? 1'b1 : 1'b0;
  /* spi_rxtx.vhdl:221:27  */
  assign n26680_o = next_cmd & cmd_valid_i;
  /* spi_rxtx.vhdl:225:29  */
  assign n26681_o = ~cmd_valid_i;
  /* spi_rxtx.vhdl:225:25  */
  assign n26682_o = next_cmd & n26681_o;
  /* spi_rxtx.vhdl:234:35  */
  assign n26685_o = state == 1'b0;
  /* spi_rxtx.vhdl:234:24  */
  assign n26686_o = n26685_o ? 1'b1 : 1'b0;
  /* spi_rxtx.vhdl:249:17  */
  assign n26691_o = end_cmd ? 1'b0 : state;
  /* spi_rxtx.vhdl:246:17  */
  assign n26692_o = start_cmd ? cmd_mode_i : cmd_mode;
  /* spi_rxtx.vhdl:246:17  */
  assign n26694_o = start_cmd ? 1'b1 : n26691_o;
  /* spi_rxtx.vhdl:240:13  */
  assign n26696_o = rst ? 3'b000 : n26692_o;
  /* spi_rxtx.vhdl:240:13  */
  assign n26698_o = rst ? 1'b0 : n26694_o;
  /* spi_rxtx.vhdl:266:29  */
  assign n26705_o = state != 1'b1;
  /* spi_rxtx.vhdl:269:72  */
  assign n26707_o = bit_count - 3'b001;
  /* spi_rxtx.vhdl:268:17  */
  assign n26708_o = sck_recv ? n26707_o : bit_count;
  /* spi_rxtx.vhdl:266:17  */
  assign n26710_o = n26705_o ? 3'b111 : n26708_o;
  /* spi_rxtx.vhdl:264:17  */
  assign n26711_o = start_cmd ? cmd_clks_i : n26710_o;
  /* spi_rxtx.vhdl:261:13  */
  assign n26713_o = rst ? 3'b000 : n26711_o;
  /* spi_rxtx.vhdl:144:20  */
  assign n26723_o = cmd_mode[2];
  /* spi_rxtx.vhdl:144:24  */
  assign n26724_o = ~n26723_o;
  /* spi_rxtx.vhdl:285:33  */
  assign n26725_o = oreg[6:0];
  /* spi_rxtx.vhdl:285:46  */
  assign n26727_o = {n26725_o, 1'b0};
  /* spi_rxtx.vhdl:148:20  */
  assign n26733_o = cmd_mode[2:1];
  /* spi_rxtx.vhdl:148:33  */
  assign n26735_o = n26733_o == 2'b10;
  /* spi_rxtx.vhdl:287:33  */
  assign n26736_o = oreg[5:0];
  /* spi_rxtx.vhdl:287:46  */
  assign n26738_o = {n26736_o, 2'b00};
  /* spi_rxtx.vhdl:289:33  */
  assign n26739_o = oreg[3:0];
  /* spi_rxtx.vhdl:289:46  */
  assign n26741_o = {n26739_o, 4'b0000};
  /* spi_rxtx.vhdl:286:17  */
  assign n26742_o = n26735_o ? n26738_o : n26741_o;
  /* spi_rxtx.vhdl:284:17  */
  assign n26743_o = n26724_o ? n26727_o : n26742_o;
  /* spi_rxtx.vhdl:282:13  */
  assign n26744_o = sck_send ? n26743_o : oreg;
  /* spi_rxtx.vhdl:280:13  */
  assign n26745_o = start_cmd ? cmd_txd_i : n26744_o;
  /* spi_rxtx.vhdl:296:22  */
  assign n26748_o = oreg[7];
  /* spi_rxtx.vhdl:298:26  */
  assign n26749_o = oreg[6];
  /* spi_rxtx.vhdl:301:26  */
  assign n26750_o = oreg[5];
  /* spi_rxtx.vhdl:302:26  */
  assign n26751_o = oreg[4];
  /* spi_rxtx.vhdl:310:22  */
  assign n26755_o = state == 1'b1;
  /* spi_rxtx.vhdl:152:20  */
  assign n26761_o = cmd_mode[2:1];
  /* spi_rxtx.vhdl:152:33  */
  assign n26763_o = n26761_o == 2'b11;
  /* spi_rxtx.vhdl:321:26  */
  assign n26765_o = 1'b1 & n26763_o;
  /* spi_rxtx.vhdl:156:20  */
  assign n26771_o = cmd_mode[0];
  /* spi_rxtx.vhdl:321:50  */
  assign n26772_o = n26765_o & n26771_o;
  /* spi_rxtx.vhdl:310:13  */
  assign n26774_o = n26775_o ? 1'b1 : 1'b0;
  /* spi_rxtx.vhdl:310:13  */
  assign n26775_o = n26755_o & n26772_o;
  /* spi_rxtx.vhdl:310:22  */
  assign n26778_o = state == 1'b1;
  /* spi_rxtx.vhdl:152:20  */
  assign n26784_o = cmd_mode[2:1];
  /* spi_rxtx.vhdl:152:33  */
  assign n26786_o = n26784_o == 2'b11;
  /* spi_rxtx.vhdl:321:26  */
  assign n26788_o = 1'b1 & n26786_o;
  /* spi_rxtx.vhdl:156:20  */
  assign n26794_o = cmd_mode[0];
  /* spi_rxtx.vhdl:321:50  */
  assign n26795_o = n26788_o & n26794_o;
  /* spi_rxtx.vhdl:310:13  */
  assign n26797_o = n26798_o ? 1'b1 : 1'b0;
  /* spi_rxtx.vhdl:310:13  */
  assign n26798_o = n26778_o & n26795_o;
  /* spi_rxtx.vhdl:310:22  */
  assign n26801_o = state == 1'b1;
  /* spi_rxtx.vhdl:148:20  */
  assign n26807_o = cmd_mode[2:1];
  /* spi_rxtx.vhdl:148:33  */
  assign n26809_o = n26807_o == 2'b10;
  /* spi_rxtx.vhdl:318:26  */
  assign n26811_o = 1'b1 & n26809_o;
  /* spi_rxtx.vhdl:156:20  */
  assign n26817_o = cmd_mode[0];
  /* spi_rxtx.vhdl:318:50  */
  assign n26818_o = n26811_o & n26817_o;
  /* spi_rxtx.vhdl:318:17  */
  assign n26820_o = n26818_o ? 1'b1 : 1'b0;
  /* spi_rxtx.vhdl:152:20  */
  assign n26826_o = cmd_mode[2:1];
  /* spi_rxtx.vhdl:152:33  */
  assign n26828_o = n26826_o == 2'b11;
  /* spi_rxtx.vhdl:321:26  */
  assign n26830_o = 1'b1 & n26828_o;
  /* spi_rxtx.vhdl:156:20  */
  assign n26836_o = cmd_mode[0];
  /* spi_rxtx.vhdl:321:50  */
  assign n26837_o = n26830_o & n26836_o;
  /* spi_rxtx.vhdl:321:17  */
  assign n26839_o = n26837_o ? 1'b1 : n26820_o;
  /* spi_rxtx.vhdl:310:13  */
  assign n26840_o = n26801_o ? n26839_o : 1'b0;
  /* spi_rxtx.vhdl:310:22  */
  assign n26843_o = state == 1'b1;
  /* spi_rxtx.vhdl:144:20  */
  assign n26849_o = cmd_mode[2];
  /* spi_rxtx.vhdl:144:24  */
  assign n26850_o = ~n26849_o;
  /* spi_rxtx.vhdl:156:20  */
  assign n26856_o = cmd_mode[0];
  /* spi_rxtx.vhdl:315:53  */
  assign n26857_o = n26850_o | n26856_o;
  /* spi_rxtx.vhdl:315:26  */
  assign n26859_o = 1'b1 & n26857_o;
  /* spi_rxtx.vhdl:310:13  */
  assign n26861_o = n26862_o ? 1'b1 : 1'b0;
  /* spi_rxtx.vhdl:310:13  */
  assign n26862_o = n26843_o & n26859_o;
  /* spi_rxtx.vhdl:354:22  */
  assign n26872_o = state == 1'b1;
  /* spi_rxtx.vhdl:354:13  */
  assign n26874_o = n26872_o ? sck_recv : 1'b0;
  /* spi_rxtx.vhdl:361:26  */
  assign n26876_o = bit_count == 3'b000;
  /* spi_rxtx.vhdl:361:34  */
  assign n26877_o = n26876_o & sck_recv;
  /* spi_rxtx.vhdl:362:42  */
  assign n26878_o = cmd_mode[0];
  /* spi_rxtx.vhdl:362:30  */
  assign n26879_o = ~n26878_o;
  /* spi_rxtx.vhdl:361:13  */
  assign n26881_o = n26877_o ? n26879_o : 1'b0;
  /* spi_rxtx.vhdl:148:20  */
  assign n26887_o = cmd_mode[2:1];
  /* spi_rxtx.vhdl:148:33  */
  assign n26889_o = n26887_o == 2'b10;
  /* spi_rxtx.vhdl:376:37  */
  assign n26890_o = ireg[5:0];
  /* spi_rxtx.vhdl:376:59  */
  assign n26891_o = dat_i_l[1];
  /* spi_rxtx.vhdl:376:50  */
  assign n26892_o = {n26890_o, n26891_o};
  /* spi_rxtx.vhdl:376:72  */
  assign n26893_o = dat_i_l[0];
  /* spi_rxtx.vhdl:376:63  */
  assign n26894_o = {n26892_o, n26893_o};
  /* spi_rxtx.vhdl:152:20  */
  assign n26900_o = cmd_mode[2:1];
  /* spi_rxtx.vhdl:152:33  */
  assign n26902_o = n26900_o == 2'b11;
  /* spi_rxtx.vhdl:378:37  */
  assign n26903_o = ireg[3:0];
  /* spi_rxtx.vhdl:378:59  */
  assign n26904_o = dat_i_l[3];
  /* spi_rxtx.vhdl:378:50  */
  assign n26905_o = {n26903_o, n26904_o};
  /* spi_rxtx.vhdl:378:72  */
  assign n26906_o = dat_i_l[2];
  /* spi_rxtx.vhdl:378:63  */
  assign n26907_o = {n26905_o, n26906_o};
  /* spi_rxtx.vhdl:378:85  */
  assign n26908_o = dat_i_l[1];
  /* spi_rxtx.vhdl:378:76  */
  assign n26909_o = {n26907_o, n26908_o};
  /* spi_rxtx.vhdl:378:98  */
  assign n26910_o = dat_i_l[0];
  /* spi_rxtx.vhdl:378:89  */
  assign n26911_o = {n26909_o, n26910_o};
  /* spi_rxtx.vhdl:381:37  */
  assign n26912_o = ireg[6:0];
  /* spi_rxtx.vhdl:381:59  */
  assign n26913_o = dat_i_l[1];
  /* spi_rxtx.vhdl:381:50  */
  assign n26914_o = {n26912_o, n26913_o};
  /* spi_rxtx.vhdl:377:21  */
  assign n26915_o = n26902_o ? n26911_o : n26914_o;
  /* spi_rxtx.vhdl:375:21  */
  assign n26916_o = n26889_o ? n26894_o : n26915_o;
  /* spi_rxtx.vhdl:173:9  */
  always @(posedge clk)
    n26923_q <= n26647_o;
  /* spi_rxtx.vhdl:173:9  */
  always @(posedge clk)
    n26924_q <= n26665_o;
  /* spi_rxtx.vhdl:173:9  */
  always @(posedge clk)
    n26925_q <= n26651_o;
  /* spi_rxtx.vhdl:173:9  */
  always @(posedge clk)
    n26926_q <= n26653_o;
  /* spi_rxtx.vhdl:173:9  */
  always @(posedge clk)
    n26927_q <= n26655_o;
  /* spi_rxtx.vhdl:239:9  */
  always @(posedge clk)
    n26928_q <= n26696_o;
  /* spi_rxtx.vhdl:278:9  */
  always @(posedge clk)
    n26929_q <= n26745_o;
  /* spi_rxtx.vhdl:342:13  */
  always @(negedge clk)
    n26930_q <= sdat_i;
  /* spi_rxtx.vhdl:351:9  */
  always @(posedge clk)
    n26931_q <= n26881_o;
  /* spi_rxtx.vhdl:351:9  */
  always @(posedge clk)
    n26932_q <= n26874_o;
  initial
    n26932_q = 1'b0;
  /* spi_rxtx.vhdl:351:9  */
  assign n26933_o = sck_recv_d ? n26916_o : ireg;
  /* spi_rxtx.vhdl:351:9  */
  always @(posedge clk)
    n26934_q <= n26933_o;
  initial
    n26934_q = 8'b00000000;
  /* spi_rxtx.vhdl:260:9  */
  always @(posedge clk)
    n26935_q <= n26713_o;
  /* spi_rxtx.vhdl:239:9  */
  always @(posedge clk)
    n26936_q <= n26698_o;
  initial
    n26936_q = 1'b0;
  /* spi_rxtx.vhdl:351:9  */
  always @(posedge clk)
    n26937_q <= dat_ack_l;
  initial
    n26937_q = 1'b0;
  /* spi_rxtx.vhdl:351:9  */
  assign n26938_o = {n26751_o, n26750_o, n26749_o, n26748_o};
  assign n26939_o = {n26774_o, n26797_o, n26840_o, n26861_o};
endmodule

module core_debug_0
  (input  clk,
   input  rst,
   input  [3:0] dmi_addr,
   input  [63:0] dmi_din,
   input  dmi_req,
   input  dmi_wr,
   input  terminate,
   input  core_stopped,
   input  [63:0] nia,
   input  [63:0] msr,
   input  dbg_gpr_ack,
   input  [63:0] dbg_gpr_data,
   input  [255:0] log_data,
   input  [31:0] log_read_addr,
   output [63:0] dmi_dout,
   output dmi_ack,
   output core_stop,
   output core_rst,
   output icache_rst,
   output dbg_gpr_req,
   output [6:0] dbg_gpr_addr,
   output [63:0] log_read_data,
   output [31:0] log_write_addr,
   output terminated_out);
  wire dmi_req_1;
  wire [63:0] stat_reg;
  wire stopping;
  wire do_step;
  wire do_reset;
  wire do_icreset;
  wire terminated;
  wire [6:0] gspr_index;
  reg [31:0] log_dmi_addr;
  reg [63:0] log_dmi_data;
  reg [63:0] log_dmi_trigger;
  reg do_log_trigger;
  wire dmi_read_log_data;
  wire dmi_read_log_data_1;
  reg [7:0] log_trigger_delay;
  wire n26304_o;
  wire n26305_o;
  wire n26307_o;
  wire n26308_o;
  wire [3:0] n26371_o;
  wire [3:0] n26372_o;
  wire [3:0] n26373_o;
  wire [3:0] n26374_o;
  wire [3:0] n26375_o;
  wire [3:0] n26376_o;
  wire [3:0] n26377_o;
  wire [3:0] n26378_o;
  wire [3:0] n26379_o;
  wire [3:0] n26380_o;
  wire [3:0] n26381_o;
  wire [3:0] n26382_o;
  wire [3:0] n26383_o;
  wire [3:0] n26384_o;
  wire [3:0] n26385_o;
  wire [3:0] n26386_o;
  wire [15:0] n26387_o;
  wire [15:0] n26388_o;
  wire [15:0] n26389_o;
  wire [15:0] n26390_o;
  wire [63:0] n26391_o;
  wire n26393_o;
  wire n26395_o;
  wire n26397_o;
  wire n26399_o;
  wire [63:0] n26400_o;
  wire n26402_o;
  wire n26404_o;
  wire n26406_o;
  wire [6:0] n26408_o;
  reg [63:0] n26409_o;
  wire [31:0] n26412_o;
  wire n26414_o;
  wire n26415_o;
  wire [31:0] n26416_o;
  wire n26418_o;
  wire [31:0] n26420_o;
  wire [31:0] n26422_o;
  wire [7:0] n26423_o;
  wire n26424_o;
  wire n26425_o;
  wire [7:0] n26427_o;
  wire n26429_o;
  wire [7:0] n26430_o;
  wire n26431_o;
  wire n26432_o;
  wire n26434_o;
  wire n26435_o;
  wire n26438_o;
  wire n26440_o;
  wire n26441_o;
  wire n26443_o;
  wire n26444_o;
  wire n26447_o;
  wire n26449_o;
  wire n26450_o;
  wire n26453_o;
  wire n26454_o;
  wire n26456_o;
  wire n26458_o;
  wire n26460_o;
  wire [6:0] n26461_o;
  wire n26463_o;
  wire [31:0] n26464_o;
  wire n26466_o;
  wire n26467_o;
  wire [61:0] n26468_o;
  wire [63:0] n26469_o;
  wire [63:0] n26470_o;
  wire [31:0] n26471_o;
  wire n26472_o;
  wire [61:0] n26473_o;
  wire [63:0] n26474_o;
  wire [63:0] n26475_o;
  wire [6:0] n26479_o;
  wire [31:0] n26480_o;
  wire n26481_o;
  wire [61:0] n26482_o;
  wire [63:0] n26483_o;
  wire [63:0] n26484_o;
  wire n26487_o;
  wire n26489_o;
  wire n26491_o;
  wire n26493_o;
  wire n26494_o;
  wire [6:0] n26495_o;
  wire [31:0] n26496_o;
  wire n26497_o;
  wire [61:0] n26498_o;
  wire [63:0] n26499_o;
  wire [63:0] n26500_o;
  wire n26503_o;
  wire n26505_o;
  wire n26507_o;
  wire n26509_o;
  wire n26510_o;
  wire [6:0] n26511_o;
  wire [31:0] n26512_o;
  wire n26513_o;
  wire [61:0] n26514_o;
  wire [63:0] n26515_o;
  wire [63:0] n26516_o;
  wire n26519_o;
  wire n26520_o;
  wire [1:0] n26521_o;
  wire [1:0] n26523_o;
  wire [1:0] n26524_o;
  wire [1:0] n26525_o;
  wire n26529_o;
  wire n26531_o;
  wire n26533_o;
  wire n26535_o;
  wire n26536_o;
  wire n26537_o;
  wire [1:0] n26538_o;
  wire [1:0] n26539_o;
  wire [29:0] n26540_o;
  wire [29:0] n26541_o;
  wire [29:0] n26542_o;
  wire n26543_o;
  wire [61:0] n26544_o;
  wire [63:0] n26545_o;
  wire [63:0] n26546_o;
  wire n26549_o;
  wire n26550_o;
  wire n26553_o;
  wire n26555_o;
  wire n26557_o;
  wire n26558_o;
  wire n26560_o;
  wire n26562_o;
  wire n26565_o;
  wire n26568_o;
  wire n26571_o;
  wire [6:0] n26572_o;
  wire [31:0] n26573_o;
  wire [31:0] n26574_o;
  wire [63:0] n26575_o;
  wire n26579_o;
  wire n26580_o;
  wire [7:0] n26582_o;
  wire n26597_o;
  wire n26598_o;
  localparam [63:0] n26599_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  localparam [31:0] n26600_o = 32'b00000000000000000000000000000001;
  reg n26601_q;
  reg n26602_q;
  reg n26603_q;
  reg n26604_q;
  reg n26605_q;
  reg n26606_q;
  reg [6:0] n26608_q;
  reg [31:0] n26609_q;
  reg [63:0] n26610_q;
  reg n26612_q;
  reg n26613_q;
  reg [7:0] n26614_q;
  assign dmi_dout = n26409_o;
  assign dmi_ack = n26305_o;
  assign core_stop = n26598_o;
  assign core_rst = do_reset;
  assign icache_rst = do_icreset;
  assign dbg_gpr_req = n26308_o;
  assign dbg_gpr_addr = gspr_index;
  assign log_read_data = n26599_o;
  assign log_write_addr = n26600_o;
  assign terminated_out = terminated;
  /* core_debug.vhdl:55:12  */
  assign dmi_req_1 = n26601_q; // (signal)
  /* core_debug.vhdl:99:12  */
  assign stat_reg = n26391_o; // (signal)
  /* core_debug.vhdl:102:12  */
  assign stopping = n26602_q; // (signal)
  /* core_debug.vhdl:103:12  */
  assign do_step = n26603_q; // (signal)
  /* core_debug.vhdl:104:12  */
  assign do_reset = n26604_q; // (signal)
  /* core_debug.vhdl:105:12  */
  assign do_icreset = n26605_q; // (signal)
  /* core_debug.vhdl:106:12  */
  assign terminated = n26606_q; // (signal)
  /* core_debug.vhdl:108:12  */
  assign gspr_index = n26608_q; // (signal)
  /* core_debug.vhdl:110:12  */
  always @*
    log_dmi_addr = n26609_q; // (isignal)
  initial
    log_dmi_addr = 32'b00000000000000000000000000000000;
  /* core_debug.vhdl:111:12  */
  always @*
    log_dmi_data = 64'b0000000000000000000000000000000000000000000000000000000000000000; // (isignal)
  initial
    log_dmi_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* core_debug.vhdl:112:12  */
  always @*
    log_dmi_trigger = n26610_q; // (isignal)
  initial
    log_dmi_trigger = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* core_debug.vhdl:113:12  */
  always @*
    do_log_trigger = 1'b0; // (isignal)
  initial
    do_log_trigger = 1'b0;
  /* core_debug.vhdl:115:12  */
  assign dmi_read_log_data = n26612_q; // (signal)
  /* core_debug.vhdl:116:12  */
  assign dmi_read_log_data_1 = n26613_q; // (signal)
  /* core_debug.vhdl:117:12  */
  always @*
    log_trigger_delay = n26614_q; // (isignal)
  initial
    log_trigger_delay = 8'b00000000;
  /* core_debug.vhdl:121:38  */
  assign n26304_o = dmi_addr != 4'b0101;
  /* core_debug.vhdl:121:24  */
  assign n26305_o = n26304_o ? dmi_req : dbg_gpr_ack;
  /* core_debug.vhdl:123:42  */
  assign n26307_o = dmi_addr == 4'b0101;
  /* core_debug.vhdl:123:28  */
  assign n26308_o = n26307_o ? dmi_req : 1'b0;
  /* dcache.vhdl:528:23  */
  assign n26371_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n26372_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n26373_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* dcache.vhdl:527:18  */
  assign n26374_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n26375_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* dcache.vhdl:527:18  */
  assign n26376_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* dcache.vhdl:525:18  */
  assign n26377_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n26378_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* dcache.vhdl:524:14  */
  assign n26379_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* dcache.vhdl:524:14  */
  assign n26380_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n26381_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* dcache.vhdl:524:14  */
  assign n26382_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n26383_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* dcache.vhdl:508:18  */
  assign n26384_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n26385_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* dcache.vhdl:507:14  */
  assign n26386_o = {1'b0, terminated, core_stopped, stopping};
  /* dcache.vhdl:507:14  */
  assign n26387_o = {n26371_o, n26372_o, n26373_o, n26374_o};
  assign n26388_o = {n26375_o, n26376_o, n26377_o, n26378_o};
  /* dcache.vhdl:507:14  */
  assign n26389_o = {n26379_o, n26380_o, n26381_o, n26382_o};
  assign n26390_o = {n26383_o, n26384_o, n26385_o, n26386_o};
  /* dcache.vhdl:508:18  */
  assign n26391_o = {n26387_o, n26388_o, n26389_o, n26390_o};
  /* core_debug.vhdl:134:25  */
  assign n26393_o = dmi_addr == 4'b0001;
  /* core_debug.vhdl:135:25  */
  assign n26395_o = dmi_addr == 4'b0010;
  /* core_debug.vhdl:136:25  */
  assign n26397_o = dmi_addr == 4'b0011;
  /* core_debug.vhdl:137:25  */
  assign n26399_o = dmi_addr == 4'b0101;
  /* core_debug.vhdl:138:24  */
  assign n26400_o = {32'b00000000000000000000000000000001, log_dmi_addr};
  /* core_debug.vhdl:138:39  */
  assign n26402_o = dmi_addr == 4'b0110;
  /* core_debug.vhdl:139:25  */
  assign n26404_o = dmi_addr == 4'b0111;
  /* core_debug.vhdl:140:25  */
  assign n26406_o = dmi_addr == 4'b1000;
  assign n26408_o = {n26406_o, n26404_o, n26402_o, n26399_o, n26397_o, n26395_o, n26393_o};
  /* core_debug.vhdl:133:5  */
  always @*
    case (n26408_o)
      7'b1000000: n26409_o = log_dmi_trigger;
      7'b0100000: n26409_o = log_dmi_data;
      7'b0010000: n26409_o = n26400_o;
      7'b0001000: n26409_o = dbg_gpr_data;
      7'b0000100: n26409_o = msr;
      7'b0000010: n26409_o = nia;
      7'b0000001: n26409_o = stat_reg;
      default: n26409_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* core_debug.vhdl:158:62  */
  assign n26412_o = {24'b0, log_trigger_delay};  //  uext
  /* core_debug.vhdl:158:62  */
  assign n26414_o = n26412_o != 32'b00000000000000000000000000000000;
  /* core_debug.vhdl:158:41  */
  assign n26415_o = do_log_trigger | n26414_o;
  /* core_debug.vhdl:159:42  */
  assign n26416_o = {24'b0, log_trigger_delay};  //  uext
  /* core_debug.vhdl:159:42  */
  assign n26418_o = n26416_o == 32'b00000000000000000000000011111111;
  /* core_debug.vhdl:163:64  */
  assign n26420_o = {24'b0, log_trigger_delay};  //  uext
  /* core_debug.vhdl:163:64  */
  assign n26422_o = n26420_o + 32'b00000000000000000000000000000001;
  /* core_debug.vhdl:163:46  */
  assign n26423_o = n26422_o[7:0];  // trunc
  /* dcache.vhdl:558:5  */
  assign n26424_o = log_dmi_trigger[1];
  /* core_debug.vhdl:158:17  */
  assign n26425_o = n26429_o ? 1'b1 : n26424_o;
  /* core_debug.vhdl:159:21  */
  assign n26427_o = n26418_o ? 8'b00000000 : n26423_o;
  /* core_debug.vhdl:158:17  */
  assign n26429_o = n26415_o & n26418_o;
  /* core_debug.vhdl:158:17  */
  assign n26430_o = n26415_o ? n26427_o : log_trigger_delay;
  /* core_debug.vhdl:168:48  */
  assign n26431_o = ~dmi_req_1;
  /* core_debug.vhdl:168:34  */
  assign n26432_o = dmi_req & n26431_o;
  /* core_debug.vhdl:173:37  */
  assign n26434_o = dmi_addr == 4'b0000;
  /* core_debug.vhdl:174:39  */
  assign n26435_o = dmi_din[1];
  /* core_debug.vhdl:174:29  */
  assign n26438_o = n26435_o ? 1'b1 : 1'b0;
  /* core_debug.vhdl:174:29  */
  assign n26440_o = n26435_o ? 1'b0 : terminated;
  /* core_debug.vhdl:178:39  */
  assign n26441_o = dmi_din[0];
  /* core_debug.vhdl:178:29  */
  assign n26443_o = n26441_o ? 1'b1 : stopping;
  /* core_debug.vhdl:181:39  */
  assign n26444_o = dmi_din[3];
  /* core_debug.vhdl:181:29  */
  assign n26447_o = n26444_o ? 1'b1 : 1'b0;
  /* core_debug.vhdl:181:29  */
  assign n26449_o = n26444_o ? 1'b0 : n26440_o;
  /* core_debug.vhdl:185:39  */
  assign n26450_o = dmi_din[2];
  /* core_debug.vhdl:185:29  */
  assign n26453_o = n26450_o ? 1'b1 : 1'b0;
  /* core_debug.vhdl:188:39  */
  assign n26454_o = dmi_din[4];
  /* core_debug.vhdl:188:29  */
  assign n26456_o = n26454_o ? 1'b0 : n26443_o;
  /* core_debug.vhdl:188:29  */
  assign n26458_o = n26454_o ? 1'b0 : n26449_o;
  /* core_debug.vhdl:192:40  */
  assign n26460_o = dmi_addr == 4'b0100;
  /* core_debug.vhdl:193:50  */
  assign n26461_o = dmi_din[6:0];
  /* core_debug.vhdl:194:40  */
  assign n26463_o = dmi_addr == 4'b0110;
  /* core_debug.vhdl:195:52  */
  assign n26464_o = dmi_din[31:0];
  /* core_debug.vhdl:197:40  */
  assign n26466_o = dmi_addr == 4'b1000;
  assign n26467_o = log_dmi_trigger[0];
  assign n26468_o = log_dmi_trigger[63:2];
  assign n26469_o = {n26468_o, n26425_o, n26467_o};
  /* core_debug.vhdl:197:25  */
  assign n26470_o = n26466_o ? dmi_din : n26469_o;
  /* core_debug.vhdl:194:25  */
  assign n26471_o = n26463_o ? n26464_o : log_dmi_addr;
  assign n26472_o = log_dmi_trigger[0];
  assign n26473_o = log_dmi_trigger[63:2];
  assign n26474_o = {n26473_o, n26425_o, n26472_o};
  /* core_debug.vhdl:194:25  */
  assign n26475_o = n26463_o ? n26474_o : n26470_o;
  /* core_debug.vhdl:192:25  */
  assign n26479_o = n26460_o ? n26461_o : gspr_index;
  /* core_debug.vhdl:192:25  */
  assign n26480_o = n26460_o ? log_dmi_addr : n26471_o;
  assign n26481_o = log_dmi_trigger[0];
  assign n26482_o = log_dmi_trigger[63:2];
  assign n26483_o = {n26482_o, n26425_o, n26481_o};
  /* core_debug.vhdl:192:25  */
  assign n26484_o = n26460_o ? n26483_o : n26475_o;
  /* core_debug.vhdl:168:17  */
  assign n26487_o = n26529_o ? n26456_o : stopping;
  /* core_debug.vhdl:173:25  */
  assign n26489_o = n26434_o ? n26447_o : 1'b0;
  /* core_debug.vhdl:173:25  */
  assign n26491_o = n26434_o ? n26438_o : 1'b0;
  /* core_debug.vhdl:173:25  */
  assign n26493_o = n26434_o ? n26453_o : 1'b0;
  /* core_debug.vhdl:168:17  */
  assign n26494_o = n26536_o ? n26458_o : terminated;
  /* core_debug.vhdl:173:25  */
  assign n26495_o = n26434_o ? gspr_index : n26479_o;
  /* core_debug.vhdl:173:25  */
  assign n26496_o = n26434_o ? log_dmi_addr : n26480_o;
  assign n26497_o = log_dmi_trigger[0];
  assign n26498_o = log_dmi_trigger[63:2];
  assign n26499_o = {n26498_o, n26425_o, n26497_o};
  /* core_debug.vhdl:173:25  */
  assign n26500_o = n26434_o ? n26499_o : n26484_o;
  /* core_debug.vhdl:169:21  */
  assign n26503_o = dmi_wr & n26434_o;
  /* core_debug.vhdl:169:21  */
  assign n26505_o = dmi_wr ? n26489_o : 1'b0;
  /* core_debug.vhdl:169:21  */
  assign n26507_o = dmi_wr ? n26491_o : 1'b0;
  /* core_debug.vhdl:169:21  */
  assign n26509_o = dmi_wr ? n26493_o : 1'b0;
  /* core_debug.vhdl:169:21  */
  assign n26510_o = dmi_wr & n26434_o;
  /* core_debug.vhdl:168:17  */
  assign n26511_o = n26537_o ? n26495_o : gspr_index;
  /* core_debug.vhdl:169:21  */
  assign n26512_o = dmi_wr ? n26496_o : log_dmi_addr;
  assign n26513_o = log_dmi_trigger[0];
  assign n26514_o = log_dmi_trigger[63:2];
  assign n26515_o = {n26514_o, n26425_o, n26513_o};
  /* core_debug.vhdl:169:21  */
  assign n26516_o = dmi_wr ? n26500_o : n26515_o;
  /* core_debug.vhdl:204:41  */
  assign n26519_o = ~dmi_read_log_data;
  /* core_debug.vhdl:204:47  */
  assign n26520_o = n26519_o & dmi_read_log_data_1;
  /* core_debug.vhdl:207:64  */
  assign n26521_o = log_dmi_addr[1:0];
  /* core_debug.vhdl:207:93  */
  assign n26523_o = n26521_o + 2'b01;
  assign n26524_o = log_dmi_addr[1:0];
  /* core_debug.vhdl:204:17  */
  assign n26525_o = n26520_o ? n26523_o : n26524_o;
  /* core_debug.vhdl:168:17  */
  assign n26529_o = n26432_o & n26503_o;
  /* core_debug.vhdl:168:17  */
  assign n26531_o = n26432_o ? n26505_o : 1'b0;
  /* core_debug.vhdl:168:17  */
  assign n26533_o = n26432_o ? n26507_o : 1'b0;
  /* core_debug.vhdl:168:17  */
  assign n26535_o = n26432_o ? n26509_o : 1'b0;
  /* core_debug.vhdl:168:17  */
  assign n26536_o = n26432_o & n26510_o;
  /* core_debug.vhdl:168:17  */
  assign n26537_o = n26432_o & dmi_wr;
  assign n26538_o = n26512_o[1:0];
  /* core_debug.vhdl:168:17  */
  assign n26539_o = n26432_o ? n26538_o : n26525_o;
  assign n26540_o = n26512_o[31:2];
  assign n26541_o = log_dmi_addr[31:2];
  /* core_debug.vhdl:168:17  */
  assign n26542_o = n26432_o ? n26540_o : n26541_o;
  assign n26543_o = log_dmi_trigger[0];
  assign n26544_o = log_dmi_trigger[63:2];
  assign n26545_o = {n26544_o, n26425_o, n26543_o};
  /* core_debug.vhdl:168:17  */
  assign n26546_o = n26432_o ? n26516_o : n26545_o;
  /* core_debug.vhdl:211:47  */
  assign n26549_o = dmi_addr == 4'b0111;
  /* core_debug.vhdl:211:34  */
  assign n26550_o = dmi_req & n26549_o;
  /* core_debug.vhdl:211:17  */
  assign n26553_o = n26550_o ? 1'b1 : 1'b0;
  /* core_debug.vhdl:220:17  */
  assign n26555_o = terminate ? 1'b1 : n26487_o;
  /* core_debug.vhdl:220:17  */
  assign n26557_o = terminate ? 1'b1 : n26494_o;
  /* core_debug.vhdl:153:13  */
  assign n26558_o = rst ? dmi_req_1 : dmi_req;
  /* core_debug.vhdl:153:13  */
  assign n26560_o = rst ? 1'b0 : n26555_o;
  /* core_debug.vhdl:153:13  */
  assign n26562_o = rst ? 1'b0 : n26531_o;
  /* core_debug.vhdl:153:13  */
  assign n26565_o = rst ? 1'b0 : n26533_o;
  /* core_debug.vhdl:153:13  */
  assign n26568_o = rst ? 1'b0 : n26535_o;
  /* core_debug.vhdl:153:13  */
  assign n26571_o = rst ? 1'b0 : n26557_o;
  /* core_debug.vhdl:153:13  */
  assign n26572_o = rst ? gspr_index : n26511_o;
  assign n26573_o = {n26542_o, n26539_o};
  /* core_debug.vhdl:153:13  */
  assign n26574_o = rst ? log_dmi_addr : n26573_o;
  /* core_debug.vhdl:153:13  */
  assign n26575_o = rst ? log_dmi_trigger : n26546_o;
  /* core_debug.vhdl:153:13  */
  assign n26579_o = rst ? dmi_read_log_data : n26553_o;
  /* core_debug.vhdl:153:13  */
  assign n26580_o = rst ? dmi_read_log_data_1 : dmi_read_log_data;
  /* core_debug.vhdl:153:13  */
  assign n26582_o = rst ? 8'b00000000 : n26430_o;
  /* core_debug.vhdl:231:31  */
  assign n26597_o = ~do_step;
  /* core_debug.vhdl:231:27  */
  assign n26598_o = stopping & n26597_o;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26601_q <= n26558_o;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26602_q <= n26560_o;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26603_q <= n26562_o;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26604_q <= n26565_o;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26605_q <= n26568_o;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26606_q <= n26571_o;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26608_q <= n26572_o;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26609_q <= n26574_o;
  initial
    n26609_q = 32'b00000000000000000000000000000000;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26610_q <= n26575_o;
  initial
    n26610_q = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26612_q <= n26579_o;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26613_q <= n26580_o;
  /* core_debug.vhdl:146:9  */
  always @(posedge clk)
    n26614_q <= n26582_o;
  initial
    n26614_q = 8'b00000000;
endmodule

module writeback
  (input  clk,
   input  rst,
   input  e_in_valid,
   input  [2:0] e_in_instr_tag,
   input  e_in_rc,
   input  e_in_mode_32bit,
   input  e_in_write_enable,
   input  [6:0] e_in_write_reg,
   input  [63:0] e_in_write_data,
   input  e_in_write_cr_enable,
   input  [7:0] e_in_write_cr_mask,
   input  [31:0] e_in_write_cr_data,
   input  e_in_write_xerc_enable,
   input  [4:0] e_in_xerc,
   input  e_in_interrupt,
   input  [11:0] e_in_intr_vec,
   input  e_in_redirect,
   input  [3:0] e_in_redir_mode,
   input  [63:0] e_in_last_nia,
   input  [63:0] e_in_br_offset,
   input  e_in_br_last,
   input  e_in_br_taken,
   input  e_in_abs_br,
   input  [15:0] e_in_srr1,
   input  [63:0] e_in_msr,
   input  l_in_valid,
   input  [2:0] l_in_instr_tag,
   input  l_in_write_enable,
   input  [6:0] l_in_write_reg,
   input  [63:0] l_in_write_data,
   input  [4:0] l_in_xerc,
   input  l_in_rc,
   input  l_in_store_done,
   input  l_in_interrupt,
   input  [11:0] l_in_intr_vec,
   input  [63:0] l_in_srr0,
   input  [15:0] l_in_srr1,
   input  fp_in_valid,
   input  fp_in_interrupt,
   input  [2:0] fp_in_instr_tag,
   input  fp_in_write_enable,
   input  [6:0] fp_in_write_reg,
   input  [63:0] fp_in_write_data,
   input  fp_in_write_cr_enable,
   input  [7:0] fp_in_write_cr_mask,
   input  [31:0] fp_in_write_cr_data,
   input  [11:0] fp_in_intr_vec,
   input  [63:0] fp_in_srr0,
   input  [15:0] fp_in_srr1,
   output [6:0] w_out_write_reg,
   output [63:0] w_out_write_data,
   output w_out_write_enable,
   output c_out_write_cr_enable,
   output [7:0] c_out_write_cr_mask,
   output [31:0] c_out_write_cr_data,
   output c_out_write_xerc_enable,
   output [4:0] c_out_write_xerc_data,
   output f_out_redirect,
   output f_out_virt_mode,
   output f_out_priv_mode,
   output f_out_big_endian,
   output f_out_mode_32bit,
   output [63:0] f_out_redirect_nia,
   output [63:0] f_out_br_nia,
   output f_out_br_last,
   output f_out_br_taken,
   output events_instr_complete,
   output events_fp_complete,
   output flush_out,
   output interrupt_out,
   output [1:0] complete_out_tag,
   output complete_out_valid);
  wire [353:0] n25972_o;
  wire [175:0] n25973_o;
  wire [209:0] n25974_o;
  wire [6:0] n25976_o;
  wire [63:0] n25977_o;
  wire n25978_o;
  wire n25980_o;
  wire [7:0] n25981_o;
  wire [31:0] n25982_o;
  wire n25983_o;
  wire [4:0] n25984_o;
  wire n25986_o;
  wire n25987_o;
  wire n25988_o;
  wire n25989_o;
  wire n25990_o;
  wire [63:0] n25991_o;
  wire [63:0] n25992_o;
  wire n25993_o;
  wire n25994_o;
  wire n25996_o;
  wire n25997_o;
  wire [1:0] n26001_o;
  wire n26002_o;
  wire [64:0] r;
  wire [64:0] rin;
  wire [64:0] n26010_o;
  wire [64:0] n26011_o;
  wire n26038_o;
  wire [2:0] n26039_o;
  wire n26040_o;
  wire [2:0] n26041_o;
  wire n26042_o;
  wire [2:0] n26043_o;
  wire [2:0] n26045_o;
  wire [2:0] n26046_o;
  wire [2:0] n26047_o;
  wire n26049_o;
  wire n26050_o;
  wire n26051_o;
  wire n26052_o;
  wire n26053_o;
  wire n26054_o;
  wire n26055_o;
  wire n26056_o;
  wire n26058_o;
  wire [63:0] n26061_o;
  wire n26068_o;
  wire [11:0] n26069_o;
  wire [63:0] n26070_o;
  wire [15:0] n26071_o;
  wire n26072_o;
  wire [11:0] n26073_o;
  wire [63:0] n26074_o;
  wire [15:0] n26075_o;
  wire n26076_o;
  wire [11:0] n26077_o;
  wire [63:0] n26078_o;
  wire [15:0] n26079_o;
  wire [63:0] n26081_o;
  wire [11:0] n26083_o;
  wire [15:0] n26085_o;
  wire [63:0] n26086_o;
  wire [11:0] n26087_o;
  wire [15:0] n26088_o;
  wire [63:0] n26089_o;
  wire [11:0] n26090_o;
  wire [15:0] n26091_o;
  wire [32:0] n26093_o;
  wire [3:0] n26094_o;
  wire [4:0] n26095_o;
  wire [5:0] n26096_o;
  wire [15:0] n26097_o;
  wire n26098_o;
  wire [6:0] n26099_o;
  wire [63:0] n26100_o;
  wire [71:0] n26102_o;
  wire [71:0] n26104_o;
  wire n26105_o;
  wire [7:0] n26107_o;
  wire [31:0] n26108_o;
  wire [40:0] n26109_o;
  localparam [40:0] n26110_o = 41'b00000000000000000000000000000000000000000;
  wire n26112_o;
  wire [4:0] n26114_o;
  wire [5:0] n26115_o;
  wire [5:0] n26117_o;
  wire n26118_o;
  wire [6:0] n26119_o;
  wire [63:0] n26120_o;
  wire [71:0] n26122_o;
  wire [71:0] n26123_o;
  wire n26124_o;
  wire [7:0] n26126_o;
  wire [31:0] n26127_o;
  wire [40:0] n26128_o;
  wire n26130_o;
  wire [6:0] n26131_o;
  wire [63:0] n26132_o;
  wire [71:0] n26134_o;
  wire [71:0] n26135_o;
  wire n26136_o;
  wire n26139_o;
  wire [4:0] n26140_o;
  wire n26141_o;
  wire [3:0] n26145_o;
  wire [8:0] n26146_o;
  wire [8:0] n26147_o;
  wire [8:0] n26148_o;
  wire [8:0] n26149_o;
  wire [8:0] n26150_o;
  wire [8:0] n26151_o;
  wire [8:0] n26152_o;
  wire [3:0] n26153_o;
  wire [3:0] n26154_o;
  wire [3:0] n26155_o;
  wire [3:0] n26156_o;
  wire [3:0] n26157_o;
  wire [3:0] n26158_o;
  wire [27:0] n26164_o;
  wire [27:0] n26165_o;
  wire [27:0] n26166_o;
  wire [27:0] n26167_o;
  wire [27:0] n26168_o;
  wire n26171_o;
  wire n26172_o;
  wire n26173_o;
  wire [31:0] n26174_o;
  wire n26175_o;
  wire n26176_o;
  wire n26177_o;
  wire n26178_o;
  wire n26179_o;
  wire [31:0] n26180_o;
  wire n26181_o;
  wire n26182_o;
  wire n26183_o;
  wire n26184_o;
  wire n26185_o;
  wire n26186_o;
  wire n26190_o;
  wire n26191_o;
  wire n26192_o;
  wire [4:0] n26193_o;
  wire n26194_o;
  wire [3:0] n26195_o;
  wire [8:0] n26196_o;
  wire [8:0] n26197_o;
  wire [3:0] n26198_o;
  wire [71:0] n26203_o;
  wire [71:0] n26204_o;
  wire [46:0] n26205_o;
  wire [46:0] n26207_o;
  wire [64:0] n26208_o;
  wire [64:0] n26209_o;
  wire [11:0] n26215_o;
  wire [71:0] n26217_o;
  wire [71:0] n26218_o;
  wire [46:0] n26221_o;
  wire n26225_o;
  wire n26227_o;
  wire n26228_o;
  wire [63:0] n26229_o;
  wire [63:0] n26230_o;
  wire [63:0] n26231_o;
  wire [11:0] n26238_o;
  wire n26241_o;
  wire [63:0] n26244_o;
  wire n26247_o;
  wire n26249_o;
  wire [30:0] n26252_o;
  wire [63:0] n26253_o;
  wire n26258_o;
  wire [63:0] n26259_o;
  wire [63:0] n26260_o;
  wire [63:0] n26261_o;
  wire [63:0] n26262_o;
  wire [63:0] n26263_o;
  wire n26264_o;
  wire n26265_o;
  wire n26266_o;
  wire n26267_o;
  wire [67:0] n26268_o;
  wire [68:0] n26269_o;
  wire n26270_o;
  wire n26271_o;
  wire [67:0] n26272_o;
  wire [67:0] n26273_o;
  wire n26274_o;
  wire [134:0] n26275_o;
  wire n26276_o;
  wire [64:0] n26277_o;
  reg [64:0] n26286_q;
  wire [1:0] n26287_o;
  assign w_out_write_reg = n25976_o;
  assign w_out_write_data = n25977_o;
  assign w_out_write_enable = n25978_o;
  assign c_out_write_cr_enable = n25980_o;
  assign c_out_write_cr_mask = n25981_o;
  assign c_out_write_cr_data = n25982_o;
  assign c_out_write_xerc_enable = n25983_o;
  assign c_out_write_xerc_data = n25984_o;
  assign f_out_redirect = n25986_o;
  assign f_out_virt_mode = n25987_o;
  assign f_out_priv_mode = n25988_o;
  assign f_out_big_endian = n25989_o;
  assign f_out_mode_32bit = n25990_o;
  assign f_out_redirect_nia = n25991_o;
  assign f_out_br_nia = n25992_o;
  assign f_out_br_last = n25993_o;
  assign f_out_br_taken = n25994_o;
  assign events_instr_complete = n25996_o;
  assign events_fp_complete = n25997_o;
  assign flush_out = n26276_o;
  assign interrupt_out = n26225_o;
  assign complete_out_tag = n26001_o;
  assign complete_out_valid = n26002_o;
  /* dcache.vhdl:1506:29  */
  assign n25972_o = {e_in_msr, e_in_srr1, e_in_abs_br, e_in_br_taken, e_in_br_last, e_in_br_offset, e_in_last_nia, e_in_redir_mode, e_in_redirect, e_in_intr_vec, e_in_interrupt, e_in_xerc, e_in_write_xerc_enable, e_in_write_cr_data, e_in_write_cr_mask, e_in_write_cr_enable, e_in_write_data, e_in_write_reg, e_in_write_enable, e_in_mode_32bit, e_in_rc, e_in_instr_tag, e_in_valid};
  /* dcache.vhdl:443:16  */
  assign n25973_o = {l_in_srr1, l_in_srr0, l_in_intr_vec, l_in_interrupt, l_in_store_done, l_in_rc, l_in_xerc, l_in_write_data, l_in_write_reg, l_in_write_enable, l_in_instr_tag, l_in_valid};
  /* dcache.vhdl:441:14  */
  assign n25974_o = {fp_in_srr1, fp_in_srr0, fp_in_intr_vec, fp_in_write_cr_data, fp_in_write_cr_mask, fp_in_write_cr_enable, fp_in_write_data, fp_in_write_reg, fp_in_write_enable, fp_in_instr_tag, fp_in_interrupt, fp_in_valid};
  assign n25976_o = n26218_o[6:0];
  /* dcache.vhdl:441:14  */
  assign n25977_o = n26218_o[70:7];
  /* dcache.vhdl:443:16  */
  assign n25978_o = n26218_o[71];
  /* dcache.vhdl:441:14  */
  assign n25980_o = n26221_o[0];
  assign n25981_o = n26221_o[8:1];
  /* dcache.vhdl:441:14  */
  assign n25982_o = n26221_o[40:9];
  /* dcache.vhdl:437:16  */
  assign n25983_o = n26221_o[41];
  /* dcache.vhdl:435:14  */
  assign n25984_o = n26221_o[46:42];
  assign n25986_o = n26275_o[0];
  /* dcache.vhdl:435:14  */
  assign n25987_o = n26275_o[1];
  /* wishbone_types.vhdl:18:14  */
  assign n25988_o = n26275_o[2];
  /* wishbone_types.vhdl:18:14  */
  assign n25989_o = n26275_o[3];
  assign n25990_o = n26275_o[4];
  /* wishbone_types.vhdl:18:14  */
  assign n25991_o = n26275_o[68:5];
  /* dcache.vhdl:1346:17  */
  assign n25992_o = n26275_o[132:69];
  assign n25993_o = n26275_o[133];
  /* dcache.vhdl:1373:21  */
  assign n25994_o = n26275_o[134];
  assign n25996_o = n26287_o[0];
  /* dcache.vhdl:501:14  */
  assign n25997_o = n26287_o[1];
  /* dcache.vhdl:1281:5  */
  assign n26001_o = n26047_o[1:0];
  /* dcache.vhdl:1284:18  */
  assign n26002_o = n26047_o[2];
  /* writeback.vhdl:39:12  */
  assign r = n26286_q; // (signal)
  /* writeback.vhdl:39:15  */
  assign rin = n26277_o; // (signal)
  assign n26010_o = {64'b0000000000000000000000000000000000000000000000000000000000000000, 1'b0};
  /* writeback.vhdl:48:13  */
  assign n26011_o = rst ? n26010_o : rin;
  /* writeback.vhdl:99:17  */
  assign n26038_o = n25972_o[0];
  /* writeback.vhdl:100:34  */
  assign n26039_o = n25972_o[3:1];
  /* writeback.vhdl:101:20  */
  assign n26040_o = n25973_o[0];
  /* writeback.vhdl:102:34  */
  assign n26041_o = n25973_o[3:1];
  /* writeback.vhdl:103:21  */
  assign n26042_o = n25974_o[0];
  /* writeback.vhdl:104:35  */
  assign n26043_o = n25974_o[4:2];
  /* writeback.vhdl:103:9  */
  assign n26045_o = n26042_o ? n26043_o : 3'b000;
  /* writeback.vhdl:101:9  */
  assign n26046_o = n26040_o ? n26041_o : n26045_o;
  /* writeback.vhdl:99:9  */
  assign n26047_o = n26038_o ? n26039_o : n26046_o;
  /* writeback.vhdl:106:47  */
  assign n26049_o = n26047_o[2];
  /* writeback.vhdl:107:37  */
  assign n26050_o = n25974_o[0];
  /* writeback.vhdl:109:22  */
  assign n26051_o = n25972_o[125];
  /* writeback.vhdl:109:40  */
  assign n26052_o = n25973_o[83];
  /* writeback.vhdl:109:32  */
  assign n26053_o = n26051_o | n26052_o;
  /* writeback.vhdl:109:59  */
  assign n26054_o = n25974_o[1];
  /* writeback.vhdl:109:50  */
  assign n26055_o = n26053_o | n26054_o;
  /* writeback.vhdl:111:14  */
  assign n26056_o = r[0];
  /* writeback.vhdl:111:20  */
  assign n26058_o = n26056_o == 1'b1;
  /* writeback.vhdl:113:35  */
  assign n26061_o = r[64:1];
  /* writeback.vhdl:123:21  */
  assign n26068_o = n25972_o[125];
  /* writeback.vhdl:124:29  */
  assign n26069_o = n25972_o[137:126];
  /* writeback.vhdl:125:42  */
  assign n26070_o = n25972_o[206:143];
  /* writeback.vhdl:126:30  */
  assign n26071_o = n25972_o[289:274];
  /* writeback.vhdl:127:24  */
  assign n26072_o = n25973_o[83];
  /* writeback.vhdl:128:29  */
  assign n26073_o = n25973_o[95:84];
  /* writeback.vhdl:129:42  */
  assign n26074_o = n25973_o[159:96];
  /* writeback.vhdl:130:30  */
  assign n26075_o = n25973_o[175:160];
  /* writeback.vhdl:131:25  */
  assign n26076_o = n25974_o[1];
  /* writeback.vhdl:132:30  */
  assign n26077_o = n25974_o[129:118];
  /* writeback.vhdl:133:43  */
  assign n26078_o = n25974_o[193:130];
  /* writeback.vhdl:134:31  */
  assign n26079_o = n25974_o[209:194];
  /* writeback.vhdl:131:13  */
  assign n26081_o = n26076_o ? n26078_o : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* writeback.vhdl:131:13  */
  assign n26083_o = n26076_o ? n26077_o : 12'b000000000000;
  /* writeback.vhdl:131:13  */
  assign n26085_o = n26076_o ? n26079_o : 16'b0000000000000000;
  /* writeback.vhdl:127:13  */
  assign n26086_o = n26072_o ? n26074_o : n26081_o;
  /* writeback.vhdl:127:13  */
  assign n26087_o = n26072_o ? n26073_o : n26083_o;
  /* writeback.vhdl:127:13  */
  assign n26088_o = n26072_o ? n26075_o : n26085_o;
  /* writeback.vhdl:123:13  */
  assign n26089_o = n26068_o ? n26070_o : n26086_o;
  /* writeback.vhdl:123:13  */
  assign n26090_o = n26068_o ? n26069_o : n26087_o;
  /* writeback.vhdl:123:13  */
  assign n26091_o = n26068_o ? n26071_o : n26088_o;
  /* writeback.vhdl:136:45  */
  assign n26093_o = n25972_o[353:321];
  /* writeback.vhdl:137:41  */
  assign n26094_o = n26091_o[14:11];
  /* writeback.vhdl:138:45  */
  assign n26095_o = n25972_o[316:312];
  /* writeback.vhdl:139:41  */
  assign n26096_o = n26091_o[5:0];
  /* writeback.vhdl:140:44  */
  assign n26097_o = n25972_o[305:290];
  /* writeback.vhdl:143:21  */
  assign n26098_o = n25972_o[6];
  /* writeback.vhdl:144:41  */
  assign n26099_o = n25972_o[13:7];
  /* writeback.vhdl:145:42  */
  assign n26100_o = n25972_o[77:14];
  assign n26102_o = {1'b1, n26100_o, n26099_o};
  /* writeback.vhdl:143:13  */
  assign n26104_o = n26098_o ? n26102_o : 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
  /* writeback.vhdl:149:21  */
  assign n26105_o = n25972_o[78];
  /* writeback.vhdl:151:45  */
  assign n26107_o = n25972_o[86:79];
  /* writeback.vhdl:152:45  */
  assign n26108_o = n25972_o[118:87];
  assign n26109_o = {n26108_o, n26107_o, 1'b1};
  /* writeback.vhdl:155:21  */
  assign n26112_o = n25972_o[119];
  /* writeback.vhdl:157:47  */
  assign n26114_o = n25972_o[124:120];
  /* dcache.vhdl:501:14  */
  assign n26115_o = {n26114_o, 1'b1};
  /* writeback.vhdl:155:13  */
  assign n26117_o = n26112_o ? n26115_o : 6'b000000;
  /* writeback.vhdl:160:22  */
  assign n26118_o = n25974_o[5];
  /* writeback.vhdl:161:42  */
  assign n26119_o = n25974_o[12:6];
  /* writeback.vhdl:162:43  */
  assign n26120_o = n25974_o[76:13];
  /* dcache.vhdl:495:14  */
  assign n26122_o = {1'b1, n26120_o, n26119_o};
  /* writeback.vhdl:160:13  */
  assign n26123_o = n26118_o ? n26122_o : n26104_o;
  /* writeback.vhdl:166:22  */
  assign n26124_o = n25974_o[77];
  /* writeback.vhdl:168:46  */
  assign n26126_o = n25974_o[85:78];
  /* writeback.vhdl:169:46  */
  assign n26127_o = n25974_o[117:86];
  /* dcache.vhdl:524:14  */
  assign n26128_o = {n26127_o, n26126_o, 1'b1};
  /* writeback.vhdl:172:21  */
  assign n26130_o = n25973_o[4];
  /* writeback.vhdl:173:41  */
  assign n26131_o = n25973_o[11:5];
  /* writeback.vhdl:174:42  */
  assign n26132_o = n25973_o[75:12];
  /* dcache.vhdl:443:16  */
  assign n26134_o = {1'b1, n26132_o, n26131_o};
  /* writeback.vhdl:172:13  */
  assign n26135_o = n26130_o ? n26134_o : n26123_o;
  /* writeback.vhdl:178:21  */
  assign n26136_o = n25973_o[81];
  /* writeback.vhdl:182:32  */
  assign n26139_o = n25973_o[82];
  /* writeback.vhdl:183:32  */
  assign n26140_o = n25973_o[80:76];
  /* writeback.vhdl:183:37  */
  assign n26141_o = n26140_o[4];
  /* dcache.vhdl:820:5  */
  assign n26145_o = {1'b0, 1'b0, n26139_o, n26141_o};
  /* dcache.vhdl:836:18  */
  assign n26146_o = {8'b10000000, 1'b1};
  assign n26147_o = n26128_o[8:0];
  /* dcache.vhdl:835:18  */
  assign n26148_o = n26109_o[8:0];
  assign n26149_o = n26110_o[8:0];
  /* writeback.vhdl:149:13  */
  assign n26150_o = n26105_o ? n26148_o : n26149_o;
  /* writeback.vhdl:166:13  */
  assign n26151_o = n26124_o ? n26147_o : n26150_o;
  /* writeback.vhdl:178:13  */
  assign n26152_o = n26136_o ? n26146_o : n26151_o;
  assign n26153_o = n26128_o[40:37];
  /* dcache.vhdl:881:39  */
  assign n26154_o = n26109_o[40:37];
  assign n26155_o = n26110_o[40:37];
  /* writeback.vhdl:149:13  */
  assign n26156_o = n26105_o ? n26154_o : n26155_o;
  /* writeback.vhdl:166:13  */
  assign n26157_o = n26124_o ? n26153_o : n26156_o;
  /* writeback.vhdl:178:13  */
  assign n26158_o = n26136_o ? n26145_o : n26157_o;
  /* dcache.vhdl:827:18  */
  assign n26164_o = n26128_o[36:9];
  assign n26165_o = n26109_o[36:9];
  /* dcache.vhdl:826:18  */
  assign n26166_o = n26110_o[36:9];
  /* writeback.vhdl:149:13  */
  assign n26167_o = n26105_o ? n26165_o : n26166_o;
  /* writeback.vhdl:166:13  */
  assign n26168_o = n26124_o ? n26164_o : n26167_o;
  /* writeback.vhdl:191:21  */
  assign n26171_o = n25972_o[4];
  /* writeback.vhdl:191:39  */
  assign n26172_o = n25972_o[6];
  /* writeback.vhdl:191:30  */
  assign n26173_o = n26171_o & n26172_o;
  /* writeback.vhdl:192:48  */
  assign n26174_o = n25972_o[45:14];
  /* writeback.vhdl:192:30  */
  assign n26175_o = |(n26174_o);
  /* writeback.vhdl:192:25  */
  assign n26176_o = ~n26175_o;
  /* writeback.vhdl:193:25  */
  assign n26177_o = n25972_o[5];
  /* writeback.vhdl:193:36  */
  assign n26178_o = ~n26177_o;
  /* writeback.vhdl:194:44  */
  assign n26179_o = n25972_o[77];
  /* writeback.vhdl:195:61  */
  assign n26180_o = n25972_o[77:46];
  /* writeback.vhdl:195:43  */
  assign n26181_o = |(n26180_o);
  /* writeback.vhdl:195:38  */
  assign n26182_o = ~n26181_o;
  /* writeback.vhdl:195:34  */
  assign n26183_o = n26176_o & n26182_o;
  /* writeback.vhdl:197:44  */
  assign n26184_o = n25972_o[45];
  /* writeback.vhdl:193:17  */
  assign n26185_o = n26178_o ? n26183_o : n26176_o;
  /* writeback.vhdl:193:17  */
  assign n26186_o = n26178_o ? n26179_o : n26184_o;
  /* writeback.vhdl:202:26  */
  assign n26190_o = ~n26186_o;
  /* writeback.vhdl:202:39  */
  assign n26191_o = ~n26185_o;
  /* writeback.vhdl:202:35  */
  assign n26192_o = n26190_o & n26191_o;
  /* writeback.vhdl:204:31  */
  assign n26193_o = n25972_o[124:120];
  /* writeback.vhdl:204:36  */
  assign n26194_o = n26193_o[4];
  /* dcache.vhdl:435:14  */
  assign n26195_o = {n26186_o, n26192_o, n26185_o, n26194_o};
  /* common.vhdl:163:14  */
  assign n26196_o = {8'b10000000, 1'b1};
  /* writeback.vhdl:191:13  */
  assign n26197_o = n26173_o ? n26196_o : n26152_o;
  /* writeback.vhdl:191:13  */
  assign n26198_o = n26173_o ? n26195_o : n26158_o;
  /* wishbone_types.vhdl:19:14  */
  assign n26203_o = {1'b1, n26089_o, 7'b0100010};
  /* writeback.vhdl:118:9  */
  assign n26204_o = n26055_o ? n26203_o : n26135_o;
  /* wishbone_types.vhdl:19:14  */
  assign n26205_o = {n26117_o, n26198_o, n26168_o, n26197_o};
  /* writeback.vhdl:118:9  */
  assign n26207_o = n26055_o ? 47'b00000000000000000000000000000000000000000000000 : n26205_o;
  assign n26208_o = {n26093_o, n26094_o, n26095_o, n26096_o, n26097_o, 1'b1};
  /* writeback.vhdl:118:9  */
  assign n26209_o = n26055_o ? n26208_o : r;
  /* writeback.vhdl:118:9  */
  assign n26215_o = n26055_o ? n26090_o : 12'b000000000000;
  /* dcache.vhdl:435:14  */
  assign n26217_o = {1'b1, n26061_o, 7'b0100011};
  /* writeback.vhdl:111:9  */
  assign n26218_o = n26058_o ? n26217_o : n26204_o;
  /* writeback.vhdl:111:9  */
  assign n26221_o = n26058_o ? 47'b00000000000000000000000000000000000000000000000 : n26207_o;
  /* writeback.vhdl:111:9  */
  assign n26225_o = n26058_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:719:9  */
  assign n26227_o = n26209_o[0];
  /* writeback.vhdl:111:9  */
  assign n26228_o = n26058_o ? 1'b0 : n26227_o;
  /* dcache.vhdl:719:9  */
  assign n26229_o = n26209_o[64:1];
  /* dcache.vhdl:719:9  */
  assign n26230_o = r[64:1];
  /* writeback.vhdl:111:9  */
  assign n26231_o = n26058_o ? n26230_o : n26229_o;
  /* writeback.vhdl:111:9  */
  assign n26238_o = n26058_o ? 12'b000000000000 : n26215_o;
  /* writeback.vhdl:210:28  */
  assign n26241_o = n25972_o[138];
  /* writeback.vhdl:211:26  */
  assign n26244_o = n25972_o[206:143];
  /* writeback.vhdl:212:27  */
  assign n26247_o = n25972_o[271];
  /* writeback.vhdl:213:28  */
  assign n26249_o = n25972_o[272];
  /* writeback.vhdl:217:61  */
  assign n26252_o = {19'b0, n26238_o};  //  uext
  /* writeback.vhdl:217:49  */
  assign n26253_o = {33'b0, n26252_o};  //  uext
  /* writeback.vhdl:224:21  */
  assign n26258_o = n25972_o[273];
  /* writeback.vhdl:225:40  */
  assign n26259_o = n25972_o[270:207];
  /* writeback.vhdl:227:67  */
  assign n26260_o = n25972_o[206:143];
  /* writeback.vhdl:227:93  */
  assign n26261_o = n25972_o[270:207];
  /* writeback.vhdl:227:77  */
  assign n26262_o = n26260_o + n26261_o;
  /* writeback.vhdl:224:13  */
  assign n26263_o = n26258_o ? n26259_o : n26262_o;
  /* writeback.vhdl:230:43  */
  assign n26264_o = n25972_o[142];
  /* writeback.vhdl:231:43  */
  assign n26265_o = n25972_o[141];
  /* writeback.vhdl:232:44  */
  assign n26266_o = n25972_o[140];
  /* writeback.vhdl:233:44  */
  assign n26267_o = n25972_o[139];
  /* dcache.vhdl:736:33  */
  assign n26268_o = {n26263_o, n26267_o, n26266_o, n26265_o, n26264_o};
  /* dcache.vhdl:711:5  */
  assign n26269_o = {n26253_o, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1};
  /* dcache.vhdl:717:18  */
  assign n26270_o = n26269_o[0];
  /* writeback.vhdl:214:9  */
  assign n26271_o = n26055_o ? n26270_o : n26241_o;
  /* dcache.vhdl:716:18  */
  assign n26272_o = n26269_o[68:1];
  /* writeback.vhdl:214:9  */
  assign n26273_o = n26055_o ? n26272_o : n26268_o;
  /* writeback.vhdl:214:9  */
  assign n26274_o = n26055_o ? 1'b0 : n26247_o;
  assign n26275_o = {n26249_o, n26274_o, n26244_o, n26273_o, n26271_o};
  /* writeback.vhdl:237:28  */
  assign n26276_o = n26275_o[0];
  assign n26277_o = {n26231_o, n26228_o};
  /* writeback.vhdl:47:9  */
  always @(posedge clk)
    n26286_q <= n26011_o;
  /* writeback.vhdl:47:9  */
  assign n26287_o = {n26050_o, n26049_o};
endmodule

module dcache_64_4_1_2_2_12_0
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  clk,
   input  rst,
   input  d_in_valid,
   input  d_in_hold,
   input  d_in_load,
   input  d_in_dcbz,
   input  d_in_nc,
   input  d_in_reserve,
   input  d_in_atomic,
   input  d_in_atomic_last,
   input  d_in_virt_mode,
   input  d_in_priv_mode,
   input  [63:0] d_in_addr,
   input  [63:0] d_in_data,
   input  [7:0] d_in_byte_sel,
   input  m_in_valid,
   input  m_in_tlbie,
   input  m_in_doall,
   input  m_in_tlbld,
   input  [63:0] m_in_addr,
   input  [63:0] m_in_pte,
   input  [28:0] snoop_in_adr,
   input  [63:0] snoop_in_dat,
   input  [7:0] snoop_in_sel,
   input  snoop_in_cyc,
   input  snoop_in_stb,
   input  snoop_in_we,
   input  [63:0] wishbone_in_dat,
   input  wishbone_in_ack,
   input  wishbone_in_stall,
   output d_out_valid,
   output [63:0] d_out_data,
   output d_out_store_done,
   output d_out_error,
   output d_out_cache_paradox,
   output m_out_stall,
   output m_out_done,
   output m_out_err,
   output [63:0] m_out_data,
   output stall_out,
   output [28:0] wishbone_out_adr,
   output [63:0] wishbone_out_dat,
   output [7:0] wishbone_out_sel,
   output wishbone_out_cyc,
   output wishbone_out_stb,
   output wishbone_out_we,
   output events_load_miss,
   output events_store_miss,
   output events_dcache_refill,
   output events_dtlb_miss,
   output events_dtlb_miss_resolved,
   output [19:0] log_out);
  wire [145:0] n23725_o;
  wire n23727_o;
  wire [63:0] n23728_o;
  wire n23729_o;
  wire n23730_o;
  wire n23731_o;
  wire [131:0] n23732_o;
  wire n23734_o;
  wire n23735_o;
  wire n23736_o;
  wire [63:0] n23737_o;
  wire [103:0] n23738_o;
  wire [28:0] n23741_o;
  wire [63:0] n23742_o;
  wire [7:0] n23743_o;
  wire n23744_o;
  wire n23745_o;
  wire n23746_o;
  wire [65:0] n23747_o;
  wire n23749_o;
  wire n23750_o;
  wire n23751_o;
  wire n23752_o;
  wire n23753_o;
  wire [47:0] cache_tag_set;
  wire [3:0] cache_valids;
  wire [3:0] dtlb_valids;
  wire [150:0] r0;
  wire r0_full;
  wire [520:0] r1;
  wire [4:0] ev;
  wire [58:0] reservation;
  wire [1:0] req_index;
  wire [4:0] req_row;
  wire [2:0] req_op;
  wire req_same_tag;
  wire req_go;
  wire [4:0] early_req_row;
  wire cancel_store;
  wire set_rsrv;
  wire clear_rsrv;
  wire r0_valid;
  wire r0_stall;
  wire use_forward_st;
  wire use_forward_rl;
  wire use_forward2;
  wire [63:0] cache_out;
  wire [63:0] ram_wr_data;
  wire [7:0] ram_wr_select;
  wire [101:0] tlb_tag_way;
  wire [127:0] tlb_pte_way;
  wire [1:0] tlb_valid_way;
  wire tlb_req_index;
  wire tlb_hit;
  wire tlb_hit_way;
  wire [63:0] pte;
  wire [55:0] ra;
  wire valid_ra;
  wire [5:0] perm_attr;
  wire rc_ok;
  wire perm_ok;
  wire access_ok;
  wire tlb_miss;
  wire [1:0] tlb_plru_victim;
  wire [47:0] snoop_tag_set;
  wire snoop_valid;
  wire [47:0] snoop_wrtag;
  wire [1:0] snoop_index;
  reg [150:0] stage_0_r;
  wire n23761_o;
  wire n23763_o;
  wire n23764_o;
  wire n23765_o;
  wire n23766_o;
  wire [63:0] n23772_o;
  wire [63:0] n23773_o;
  wire n23775_o;
  wire n23776_o;
  wire n23777_o;
  wire [7:0] n23781_o;
  wire [73:0] n23782_o;
  wire [150:0] n23788_o;
  wire [3:0] n23789_o;
  wire [142:0] n23790_o;
  wire n23791_o;
  wire n23792_o;
  wire n23793_o;
  wire n23794_o;
  wire n23795_o;
  wire [3:0] n23796_o;
  wire [3:0] n23797_o;
  wire [1:0] n23798_o;
  wire [1:0] n23799_o;
  wire [1:0] n23800_o;
  wire [142:0] n23801_o;
  wire [142:0] n23802_o;
  wire n23803_o;
  wire n23804_o;
  wire n23805_o;
  wire n23806_o;
  wire n23807_o;
  wire n23808_o;
  wire n23809_o;
  wire [150:0] n23810_o;
  wire [150:0] n23811_o;
  wire [145:0] n23812_o;
  wire n23813_o;
  wire n23814_o;
  wire n23815_o;
  wire [63:0] n23816_o;
  wire [145:0] n23817_o;
  wire n23818_o;
  wire [63:0] n23819_o;
  wire [63:0] n23820_o;
  wire n23821_o;
  wire n23822_o;
  wire [73:0] n23823_o;
  wire [73:0] n23824_o;
  wire [73:0] n23825_o;
  wire [63:0] n23826_o;
  wire [63:0] n23827_o;
  wire [11:0] n23828_o;
  wire [11:0] n23829_o;
  wire [11:0] n23830_o;
  wire n23831_o;
  wire n23832_o;
  wire n23833_o;
  wire [150:0] n23834_o;
  wire [150:0] n23835_o;
  wire n23837_o;
  wire [150:0] n23840_o;
  reg [150:0] n23843_q;
  wire n23845_o;
  wire n23846_o;
  wire n23847_o;
  wire n23848_o;
  wire n23849_o;
  wire n23850_o;
  wire n23851_o;
  wire n23852_o;
  wire n23853_o;
  wire n23854_o;
  wire n23859_o;
  wire n23860_o;
  wire n23861_o;
  wire n23862_o;
  wire n23864_o;
  wire n23866_o;
  wire maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_acc;
  wire maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_acc_en;
  wire maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_out;
  wire maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_lru;
  wire n23889_o;
  wire [31:0] n23890_o;
  wire n23892_o;
  wire n23893_o;
  wire n23895_o;
  wire n23896_o;
  wire maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_acc;
  wire maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_acc_en;
  wire maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_out;
  wire maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_lru;
  wire n23902_o;
  wire [31:0] n23903_o;
  wire n23905_o;
  wire n23906_o;
  wire n23908_o;
  wire n23909_o;
  wire n23916_o;
  wire [50:0] n23918_o;
  wire n23919_o;
  wire [50:0] n23926_o;
  wire n23927_o;
  wire n23928_o;
  wire n23931_o;
  wire n23933_o;
  wire [50:0] n23940_o;
  wire n23941_o;
  wire n23942_o;
  wire n23945_o;
  wire n23948_o;
  wire n23949_o;
  wire [63:0] n23967_o;
  wire [145:0] n23968_o;
  wire n23969_o;
  wire n23970_o;
  wire n23971_o;
  wire [145:0] n23972_o;
  wire n23973_o;
  wire n23974_o;
  wire n23975_o;
  wire n23976_o;
  wire [145:0] n23977_o;
  wire n23978_o;
  wire [43:0] n23979_o;
  wire [8:0] n23980_o;
  wire [52:0] n23981_o;
  wire [55:0] n23983_o;
  wire n23990_o;
  wire n23993_o;
  wire n23995_o;
  wire n23997_o;
  wire n23999_o;
  wire n24001_o;
  wire [5:0] n24002_o;
  wire [52:0] n24003_o;
  wire [55:0] n24005_o;
  wire [55:0] n24006_o;
  wire [5:0] n24008_o;
  wire n24019_o;
  wire n24020_o;
  wire n24021_o;
  wire n24022_o;
  wire n24023_o;
  wire n24024_o;
  wire n24025_o;
  wire n24029_o;
  wire [3:0] n24035_o;
  wire n24037_o;
  wire n24041_o;
  wire [50:0] n24042_o;
  wire [145:0] n24062_o;
  wire [63:0] n24063_o;
  wire n24082_o;
  wire [3:0] n24088_o;
  wire [3:0] n24095_o;
  wire [3:0] n24102_o;
  wire [3:0] n24103_o;
  wire n24129_o;
  wire [63:0] n24131_o;
  wire [1:0] n24136_o;
  wire [63:0] n24139_o;
  wire [1:0] n24144_o;
  wire [1:0] n24146_o;
  wire [1:0] n24147_o;
  wire [28:0] n24160_o;
  localparam [63:0] n24166_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] n24167_o;
  wire [2:0] n24168_o;
  wire [63:0] n24169_o;
  wire [55:0] n24174_o;
  wire [1:0] n24180_o;
  wire [47:0] n24191_o;
  wire [1:0] n24197_o;
  wire [103:0] n24199_o;
  wire n24200_o;
  wire n24201_o;
  wire n24202_o;
  wire n24203_o;
  wire n24204_o;
  wire n24205_o;
  wire n24206_o;
  wire n24207_o;
  wire n24208_o;
  wire n24209_o;
  wire n24211_o;
  wire [145:0] n24237_o;
  wire [63:0] n24238_o;
  wire [1:0] n24243_o;
  wire [145:0] n24246_o;
  wire [63:0] n24247_o;
  wire [4:0] n24252_o;
  wire n24260_o;
  wire n24261_o;
  wire n24262_o;
  wire n24263_o;
  wire n24264_o;
  wire n24265_o;
  wire n24266_o;
  wire n24267_o;
  wire [145:0] n24268_o;
  wire n24269_o;
  wire [63:0] n24276_o;
  wire [43:0] n24277_o;
  wire [11:0] n24278_o;
  wire [55:0] n24279_o;
  wire [47:0] n24285_o;
  wire [1:0] n24287_o;
  wire n24290_o;
  wire n24296_o;
  wire n24297_o;
  wire n24298_o;
  wire n24299_o;
  wire n24302_o;
  wire [47:0] n24304_o;
  wire n24305_o;
  wire n24308_o;
  localparam [1:0] n24309_o = 2'b00;
  wire n24310_o;
  wire [47:0] n24311_o;
  wire n24312_o;
  wire n24315_o;
  localparam [1:0] n24316_o = 2'b00;
  wire n24317_o;
  wire [63:0] n24324_o;
  wire [43:0] n24325_o;
  wire [11:0] n24326_o;
  wire [55:0] n24327_o;
  wire [47:0] n24333_o;
  wire [1:0] n24335_o;
  wire n24338_o;
  wire n24344_o;
  wire n24345_o;
  wire n24346_o;
  wire n24347_o;
  wire n24350_o;
  wire [47:0] n24352_o;
  wire n24353_o;
  wire n24355_o;
  wire [47:0] n24356_o;
  wire n24357_o;
  wire n24359_o;
  wire [1:0] n24361_o;
  wire [1:0] n24367_o;
  wire [1:0] n24370_o;
  wire n24373_o;
  wire n24375_o;
  wire n24377_o;
  wire [145:0] n24379_o;
  wire [63:0] n24380_o;
  wire [47:0] n24385_o;
  wire [1:0] n24387_o;
  wire n24390_o;
  wire n24396_o;
  wire n24397_o;
  wire n24400_o;
  wire [47:0] n24401_o;
  wire n24402_o;
  wire n24405_o;
  wire [47:0] n24406_o;
  wire n24407_o;
  wire n24410_o;
  wire n24411_o;
  wire n24421_o;
  wire n24425_o;
  wire [4:0] n24427_o;
  wire [31:0] n24428_o;
  wire [31:0] n24429_o;
  wire n24430_o;
  wire n24431_o;
  wire n24432_o;
  wire [1:0] n24433_o;
  wire n24435_o;
  wire n24436_o;
  wire n24437_o;
  wire n24440_o;
  wire n24442_o;
  wire n24445_o;
  wire [4:0] n24447_o;
  wire [31:0] n24448_o;
  wire [31:0] n24449_o;
  wire n24450_o;
  wire n24451_o;
  wire n24452_o;
  wire n24454_o;
  wire [1:0] n24463_o;
  wire n24465_o;
  wire [31:0] n24466_o;
  wire [1:0] n24467_o;
  wire [31:0] n24468_o;
  wire n24469_o;
  wire n24470_o;
  wire n24471_o;
  wire [145:0] n24472_o;
  wire n24473_o;
  wire n24474_o;
  wire [31:0] n24475_o;
  wire [2:0] n24476_o;
  wire [2:0] n24479_o;
  wire n24482_o;
  wire n24483_o;
  wire n24484_o;
  wire n24485_o;
  wire [145:0] n24486_o;
  wire n24487_o;
  wire n24488_o;
  wire n24489_o;
  wire n24490_o;
  wire [145:0] n24491_o;
  wire n24492_o;
  wire n24493_o;
  wire n24494_o;
  wire n24495_o;
  wire n24496_o;
  wire [145:0] n24497_o;
  wire n24498_o;
  wire n24499_o;
  wire n24500_o;
  wire n24501_o;
  wire n24502_o;
  wire n24503_o;
  wire n24504_o;
  wire [145:0] n24505_o;
  wire n24506_o;
  wire n24507_o;
  wire n24508_o;
  wire n24509_o;
  wire [145:0] n24510_o;
  wire n24511_o;
  wire [1:0] n24512_o;
  wire [2:0] n24513_o;
  wire n24515_o;
  wire n24517_o;
  wire n24519_o;
  wire n24521_o;
  wire n24523_o;
  wire n24525_o;
  wire n24527_o;
  wire n24529_o;
  wire [7:0] n24530_o;
  reg [2:0] n24540_o;
  wire [2:0] n24542_o;
  wire [2:0] n24545_o;
  wire [2:0] n24548_o;
  wire n24551_o;
  wire n24552_o;
  wire [63:0] n24554_o;
  wire [4:0] n24559_o;
  wire [63:0] n24562_o;
  wire [4:0] n24567_o;
  wire [4:0] n24569_o;
  wire [4:0] n24570_o;
  wire [103:0] n24578_o;
  wire [145:0] n24580_o;
  wire n24581_o;
  wire n24582_o;
  wire [145:0] n24583_o;
  wire n24584_o;
  wire [145:0] n24585_o;
  wire n24586_o;
  wire [145:0] n24587_o;
  wire n24588_o;
  wire n24589_o;
  wire n24590_o;
  wire [57:0] n24591_o;
  wire [57:0] n24592_o;
  wire n24593_o;
  wire n24594_o;
  wire n24597_o;
  wire n24599_o;
  wire n24601_o;
  wire n24603_o;
  wire n24605_o;
  wire n24608_o;
  wire n24611_o;
  wire n24617_o;
  wire [57:0] n24620_o;
  wire [58:0] n24621_o;
  wire [58:0] n24622_o;
  wire n24623_o;
  wire n24624_o;
  wire [57:0] n24625_o;
  wire [57:0] n24626_o;
  wire [57:0] n24627_o;
  wire [58:0] n24628_o;
  wire [58:0] n24629_o;
  wire n24630_o;
  wire n24631_o;
  wire [57:0] n24632_o;
  wire [57:0] n24633_o;
  wire [57:0] n24634_o;
  wire [58:0] n24635_o;
  wire n24639_o;
  wire [63:0] n24640_o;
  wire n24641_o;
  wire n24642_o;
  wire n24643_o;
  wire n24644_o;
  wire n24645_o;
  wire n24646_o;
  wire [63:0] n24647_o;
  wire [134:0] n24657_o;
  wire [63:0] n24658_o;
  wire n24659_o;
  wire [63:0] n24660_o;
  wire [63:0] n24661_o;
  wire n24662_o;
  wire n24663_o;
  wire [63:0] n24664_o;
  wire [134:0] n24666_o;
  wire [7:0] n24667_o;
  wire n24668_o;
  wire [7:0] n24669_o;
  wire rams_n1_do_read;
  wire [4:0] rams_n1_rd_addr;
  wire [4:0] rams_n1_wr_addr;
  wire [7:0] rams_n1_wr_sel_m;
  wire [63:0] rams_n1_dout;
  wire [63:0] rams_n1_way_rd_data;
  wire [4:0] n24675_o;
  wire n24677_o;
  wire [1:0] n24678_o;
  wire n24680_o;
  wire n24681_o;
  wire n24682_o;
  wire n24683_o;
  wire n24685_o;
  wire [7:0] n24687_o;
  wire n24701_o;
  wire n24704_o;
  wire n24705_o;
  wire n24706_o;
  wire [1:0] n24708_o;
  wire n24709_o;
  wire n24710_o;
  wire n24711_o;
  wire n24712_o;
  wire [1:0] n24715_o;
  wire [1:0] n24717_o;
  wire [1:0] n24718_o;
  wire [7:0] n24719_o;
  wire n24721_o;
  wire [7:0] n24722_o;
  wire n24724_o;
  wire [7:0] n24725_o;
  wire n24727_o;
  wire [7:0] n24728_o;
  wire [2:0] n24729_o;
  reg [7:0] n24730_o;
  wire n24731_o;
  wire n24732_o;
  wire n24733_o;
  wire [1:0] n24735_o;
  wire n24736_o;
  wire n24737_o;
  wire n24738_o;
  wire n24739_o;
  wire [1:0] n24742_o;
  wire [1:0] n24744_o;
  wire [1:0] n24745_o;
  wire [7:0] n24746_o;
  wire n24748_o;
  wire [7:0] n24749_o;
  wire n24751_o;
  wire [7:0] n24752_o;
  wire n24754_o;
  wire [7:0] n24755_o;
  wire [2:0] n24756_o;
  reg [7:0] n24757_o;
  wire n24758_o;
  wire n24759_o;
  wire n24760_o;
  wire [1:0] n24762_o;
  wire n24763_o;
  wire n24764_o;
  wire n24765_o;
  wire n24766_o;
  wire [1:0] n24769_o;
  wire [1:0] n24771_o;
  wire [1:0] n24772_o;
  wire [7:0] n24773_o;
  wire n24775_o;
  wire [7:0] n24776_o;
  wire n24778_o;
  wire [7:0] n24779_o;
  wire n24781_o;
  wire [7:0] n24782_o;
  wire [2:0] n24783_o;
  reg [7:0] n24784_o;
  wire n24785_o;
  wire n24786_o;
  wire n24787_o;
  wire [1:0] n24789_o;
  wire n24790_o;
  wire n24791_o;
  wire n24792_o;
  wire n24793_o;
  wire [1:0] n24796_o;
  wire [1:0] n24798_o;
  wire [1:0] n24799_o;
  wire [7:0] n24800_o;
  wire n24802_o;
  wire [7:0] n24803_o;
  wire n24805_o;
  wire [7:0] n24806_o;
  wire n24808_o;
  wire [7:0] n24809_o;
  wire [2:0] n24810_o;
  reg [7:0] n24811_o;
  wire n24812_o;
  wire n24813_o;
  wire n24814_o;
  wire [1:0] n24816_o;
  wire n24817_o;
  wire n24818_o;
  wire n24819_o;
  wire n24820_o;
  wire [1:0] n24823_o;
  wire [1:0] n24825_o;
  wire [1:0] n24826_o;
  wire [7:0] n24827_o;
  wire n24829_o;
  wire [7:0] n24830_o;
  wire n24832_o;
  wire [7:0] n24833_o;
  wire n24835_o;
  wire [7:0] n24836_o;
  wire [2:0] n24837_o;
  reg [7:0] n24838_o;
  wire n24839_o;
  wire n24840_o;
  wire n24841_o;
  wire [1:0] n24843_o;
  wire n24844_o;
  wire n24845_o;
  wire n24846_o;
  wire n24847_o;
  wire [1:0] n24850_o;
  wire [1:0] n24852_o;
  wire [1:0] n24853_o;
  wire [7:0] n24854_o;
  wire n24856_o;
  wire [7:0] n24857_o;
  wire n24859_o;
  wire [7:0] n24860_o;
  wire n24862_o;
  wire [7:0] n24863_o;
  wire [2:0] n24864_o;
  reg [7:0] n24865_o;
  wire n24866_o;
  wire n24867_o;
  wire n24868_o;
  wire [1:0] n24870_o;
  wire n24871_o;
  wire n24872_o;
  wire n24873_o;
  wire n24874_o;
  wire [1:0] n24877_o;
  wire [1:0] n24879_o;
  wire [1:0] n24880_o;
  wire [7:0] n24881_o;
  wire n24883_o;
  wire [7:0] n24884_o;
  wire n24886_o;
  wire [7:0] n24887_o;
  wire n24889_o;
  wire [7:0] n24890_o;
  wire [2:0] n24891_o;
  reg [7:0] n24892_o;
  wire n24893_o;
  wire n24894_o;
  wire n24895_o;
  wire [1:0] n24897_o;
  wire n24898_o;
  wire n24899_o;
  wire n24900_o;
  wire n24901_o;
  wire [1:0] n24904_o;
  wire [1:0] n24906_o;
  wire [1:0] n24907_o;
  wire [7:0] n24908_o;
  wire n24910_o;
  wire [7:0] n24911_o;
  wire n24913_o;
  wire [7:0] n24914_o;
  wire n24916_o;
  wire [7:0] n24917_o;
  wire [2:0] n24918_o;
  reg [7:0] n24919_o;
  wire [63:0] n24920_o;
  wire [47:0] n24921_o;
  wire [4:0] n24922_o;
  wire n24923_o;
  wire [1:0] n24924_o;
  wire n24926_o;
  wire n24927_o;
  wire n24928_o;
  wire n24930_o;
  wire n24932_o;
  wire n24935_o;
  wire n24937_o;
  wire n24939_o;
  wire n24940_o;
  wire n24943_o;
  wire n24945_o;
  wire n24946_o;
  wire n24947_o;
  wire n24948_o;
  wire [1:0] n24952_o;
  wire [1:0] n24953_o;
  wire n24954_o;
  wire [1:0] n24955_o;
  wire n24957_o;
  wire n24960_o;
  wire [196:0] n24961_o;
  wire [2:0] n24962_o;
  wire n25002_o;
  wire n25003_o;
  wire n25004_o;
  wire n25005_o;
  wire n25007_o;
  wire n25009_o;
  wire n25010_o;
  wire n25011_o;
  wire n25012_o;
  wire n25015_o;
  wire n25016_o;
  wire n25017_o;
  wire n25018_o;
  wire n25024_o;
  wire n25025_o;
  wire [1:0] n25027_o;
  wire [3:0] n25031_o;
  wire n25032_o;
  wire [1:0] n25033_o;
  wire [47:0] n25037_o;
  wire n25042_o;
  wire n25043_o;
  wire n25044_o;
  wire [134:0] n25045_o;
  wire n25046_o;
  wire [145:0] n25047_o;
  wire n25048_o;
  wire [145:0] n25049_o;
  wire n25050_o;
  wire n25052_o;
  wire [145:0] n25053_o;
  wire [63:0] n25054_o;
  wire [63:0] n25055_o;
  wire [63:0] n25056_o;
  wire [63:0] n25057_o;
  wire [145:0] n25058_o;
  wire n25059_o;
  wire [145:0] n25060_o;
  wire n25061_o;
  wire [145:0] n25062_o;
  wire n25063_o;
  wire n25064_o;
  wire n25065_o;
  wire n25066_o;
  wire n25067_o;
  wire n25068_o;
  wire n25069_o;
  wire [145:0] n25071_o;
  wire [7:0] n25072_o;
  wire [7:0] n25073_o;
  wire n25075_o;
  wire n25077_o;
  wire n25078_o;
  wire n25080_o;
  wire n25081_o;
  wire n25083_o;
  wire n25084_o;
  wire [134:0] n25085_o;
  wire n25087_o;
  wire n25088_o;
  wire n25091_o;
  wire n25092_o;
  wire [134:0] n25095_o;
  wire [134:0] n25096_o;
  wire [1:0] n25097_o;
  wire [55:0] n25099_o;
  wire [28:0] n25104_o;
  wire [7:0] n25105_o;
  wire [63:0] n25106_o;
  wire n25107_o;
  wire [55:0] n25109_o;
  wire [1:0] n25114_o;
  wire [55:0] n25117_o;
  wire [4:0] n25122_o;
  wire [55:0] n25126_o;
  wire [4:0] n25131_o;
  wire [2:0] n25140_o;
  wire [2:0] n25142_o;
  wire [55:0] n25144_o;
  wire [47:0] n25149_o;
  wire [2:0] n25162_o;
  wire n25164_o;
  wire n25172_o;
  wire n25178_o;
  wire n25179_o;
  wire n25180_o;
  wire n25185_o;
  wire n25186_o;
  wire n25189_o;
  wire n25190_o;
  wire [2:0] n25191_o;
  wire n25193_o;
  wire n25195_o;
  wire [2:0] n25197_o;
  wire n25199_o;
  wire n25201_o;
  wire n25202_o;
  wire [1:0] n25203_o;
  wire n25204_o;
  wire n25205_o;
  wire n25206_o;
  wire [2:0] n25207_o;
  wire [2:0] n25208_o;
  wire n25209_o;
  wire n25210_o;
  wire [2:0] n25214_o;
  wire n25216_o;
  wire n25218_o;
  wire n25220_o;
  wire n25222_o;
  wire n25223_o;
  wire n25225_o;
  wire n25227_o;
  wire n25229_o;
  wire [6:0] n25230_o;
  reg n25232_o;
  wire [1:0] n25233_o;
  reg [1:0] n25235_o;
  reg n25237_o;
  reg n25239_o;
  reg n25241_o;
  wire n25242_o;
  reg n25244_o;
  wire n25245_o;
  reg n25247_o;
  wire n25248_o;
  reg n25250_o;
  wire [2:0] n25251_o;
  reg [2:0] n25253_o;
  reg n25255_o;
  reg n25257_o;
  reg n25259_o;
  reg n25261_o;
  wire n25263_o;
  wire n25264_o;
  wire n25265_o;
  wire [103:0] n25266_o;
  wire n25267_o;
  wire n25268_o;
  wire [103:0] n25270_o;
  wire [28:0] n25271_o;
  wire [2:0] n25272_o;
  wire [2:0] n25277_o;
  wire n25278_o;
  wire n25280_o;
  wire n25281_o;
  wire [103:0] n25283_o;
  wire [28:0] n25284_o;
  wire [2:0] n25291_o;
  wire [2:0] n25294_o;
  wire [25:0] n25296_o;
  wire [28:0] n25297_o;
  wire [28:0] n25298_o;
  wire [28:0] n25299_o;
  wire n25301_o;
  wire n25302_o;
  wire [4:0] n25303_o;
  wire [31:0] n25304_o;
  wire [2:0] n25305_o;
  wire [2:0] n25308_o;
  wire [7:0] n25310_o;
  wire n25313_o;
  wire [134:0] n25314_o;
  wire n25315_o;
  wire n25316_o;
  wire n25317_o;
  wire n25318_o;
  wire n25319_o;
  wire [134:0] n25320_o;
  wire [2:0] n25321_o;
  wire n25323_o;
  wire n25324_o;
  wire n25325_o;
  wire [4:0] n25326_o;
  wire [31:0] n25327_o;
  wire [134:0] n25329_o;
  wire [55:0] n25330_o;
  wire [4:0] n25335_o;
  wire [31:0] n25337_o;
  wire n25338_o;
  wire n25339_o;
  wire n25342_o;
  wire n25343_o;
  wire n25346_o;
  wire n25347_o;
  wire n25348_o;
  wire n25349_o;
  wire n25350_o;
  wire n25351_o;
  wire [4:0] n25353_o;
  wire [2:0] n25354_o;
  wire [2:0] n25367_o;
  wire n25368_o;
  wire [1:0] n25370_o;
  wire [1:0] n25372_o;
  wire n25376_o;
  wire n25377_o;
  wire [3:0] n25379_o;
  wire [1:0] n25380_o;
  wire [1:0] n25381_o;
  wire n25382_o;
  wire n25383_o;
  wire n25384_o;
  wire [4:0] n25386_o;
  wire [2:0] n25396_o;
  wire [2:0] n25399_o;
  wire [1:0] n25400_o;
  wire [4:0] n25401_o;
  wire n25403_o;
  wire n25404_o;
  wire n25406_o;
  wire n25407_o;
  wire n25409_o;
  wire [4:0] n25410_o;
  wire [4:0] n25411_o;
  wire [7:0] n25412_o;
  wire [7:0] n25413_o;
  wire n25414_o;
  wire n25415_o;
  wire n25416_o;
  wire n25418_o;
  wire [103:0] n25419_o;
  wire n25420_o;
  wire n25421_o;
  wire [2:0] n25422_o;
  wire n25423_o;
  wire n25424_o;
  wire n25425_o;
  wire n25426_o;
  wire [2:0] n25428_o;
  wire [2:0] n25430_o;
  wire [2:0] n25431_o;
  wire [2:0] n25432_o;
  wire n25433_o;
  wire n25434_o;
  wire n25435_o;
  wire [4:0] n25436_o;
  wire [63:0] n25437_o;
  wire [7:0] n25438_o;
  wire [71:0] n25439_o;
  wire [4:0] n25440_o;
  wire [4:0] n25441_o;
  wire [71:0] n25442_o;
  wire [71:0] n25443_o;
  wire n25445_o;
  wire n25446_o;
  wire n25447_o;
  wire n25448_o;
  wire n25449_o;
  wire n25450_o;
  wire [2:0] n25451_o;
  wire n25453_o;
  wire [2:0] n25454_o;
  wire n25456_o;
  wire n25457_o;
  wire n25458_o;
  wire [55:0] n25461_o;
  wire [4:0] n25466_o;
  wire [2:0] n25468_o;
  wire n25470_o;
  wire n25472_o;
  wire n25478_o;
  wire n25479_o;
  wire n25480_o;
  wire n25481_o;
  wire [4:0] n25482_o;
  wire [4:0] n25483_o;
  wire n25484_o;
  wire n25485_o;
  wire n25488_o;
  wire [5:0] n25489_o;
  wire n25490_o;
  wire n25491_o;
  wire [4:0] n25492_o;
  wire [5:0] n25493_o;
  wire [5:0] n25494_o;
  wire n25496_o;
  wire n25497_o;
  wire n25498_o;
  wire n25500_o;
  wire n25501_o;
  wire n25502_o;
  wire n25503_o;
  wire n25504_o;
  wire n25506_o;
  wire n25507_o;
  wire [1:0] n25511_o;
  wire [1:0] n25512_o;
  wire [1:0] n25513_o;
  wire n25514_o;
  wire [1:0] n25515_o;
  wire [1:0] n25516_o;
  wire n25519_o;
  wire n25520_o;
  wire [1:0] n25521_o;
  wire [1:0] n25522_o;
  wire n25523_o;
  wire n25525_o;
  wire n25526_o;
  wire n25527_o;
  wire n25529_o;
  wire n25530_o;
  wire n25531_o;
  wire n25535_o;
  wire n25536_o;
  wire n25539_o;
  wire n25540_o;
  wire [1:0] n25543_o;
  wire n25544_o;
  wire [1:0] n25545_o;
  wire [1:0] n25546_o;
  wire n25547_o;
  wire n25548_o;
  wire [1:0] n25549_o;
  wire [1:0] n25550_o;
  wire n25551_o;
  wire n25552_o;
  wire n25554_o;
  wire [3:0] n25555_o;
  reg [3:0] n25557_o;
  reg n25559_o;
  wire n25560_o;
  wire n25561_o;
  wire n25562_o;
  wire n25563_o;
  wire n25564_o;
  reg n25566_o;
  reg [1:0] n25568_o;
  wire n25569_o;
  reg n25571_o;
  reg n25573_o;
  reg n25575_o;
  wire n25576_o;
  reg n25578_o;
  wire [4:0] n25579_o;
  wire [4:0] n25580_o;
  wire [4:0] n25581_o;
  wire [4:0] n25582_o;
  reg [4:0] n25584_o;
  wire [23:0] n25585_o;
  wire [23:0] n25586_o;
  wire [23:0] n25587_o;
  reg [23:0] n25589_o;
  wire [63:0] n25590_o;
  wire [63:0] n25591_o;
  reg [63:0] n25593_o;
  wire [7:0] n25594_o;
  wire [7:0] n25595_o;
  reg [7:0] n25597_o;
  wire n25598_o;
  wire n25599_o;
  reg n25601_o;
  wire n25602_o;
  wire n25603_o;
  reg n25605_o;
  wire n25606_o;
  reg n25608_o;
  wire [47:0] n25609_o;
  reg [47:0] n25611_o;
  wire [4:0] n25612_o;
  reg [4:0] n25614_o;
  wire [1:0] n25615_o;
  reg [1:0] n25617_o;
  wire [2:0] n25618_o;
  reg [2:0] n25620_o;
  wire n25621_o;
  wire n25622_o;
  reg n25624_o;
  wire n25625_o;
  wire n25626_o;
  reg n25628_o;
  wire n25629_o;
  wire n25630_o;
  reg n25632_o;
  wire n25633_o;
  wire n25634_o;
  reg n25636_o;
  wire n25637_o;
  wire n25638_o;
  reg n25640_o;
  wire n25641_o;
  wire n25642_o;
  reg n25644_o;
  wire n25645_o;
  wire n25646_o;
  reg n25648_o;
  wire n25649_o;
  wire n25650_o;
  reg n25652_o;
  wire [2:0] n25653_o;
  reg [2:0] n25655_o;
  reg n25657_o;
  reg n25659_o;
  reg n25661_o;
  reg n25663_o;
  wire n25664_o;
  wire n25665_o;
  wire n25666_o;
  wire n25667_o;
  wire n25668_o;
  wire [132:0] n25669_o;
  wire [132:0] n25670_o;
  wire [132:0] n25671_o;
  wire [132:0] n25672_o;
  wire [132:0] n25673_o;
  reg n25675_o;
  reg n25677_o;
  reg n25679_o;
  wire [3:0] n25685_o;
  wire [3:0] n25686_o;
  wire [134:0] n25687_o;
  wire [181:0] n25688_o;
  wire [29:0] n25689_o;
  wire [1:0] n25690_o;
  wire n25691_o;
  wire [134:0] n25692_o;
  wire [134:0] n25693_o;
  wire [1:0] n25694_o;
  wire [1:0] n25695_o;
  wire [2:0] n25696_o;
  wire [2:0] n25697_o;
  wire [2:0] n25698_o;
  wire [29:0] n25699_o;
  wire [29:0] n25700_o;
  wire [71:0] n25701_o;
  wire [71:0] n25702_o;
  wire [71:0] n25703_o;
  wire [1:0] n25704_o;
  wire [1:0] n25705_o;
  wire [71:0] n25706_o;
  wire [71:0] n25707_o;
  wire [71:0] n25708_o;
  wire n25709_o;
  wire n25710_o;
  wire n25711_o;
  wire [2:0] n25712_o;
  wire [2:0] n25713_o;
  wire [2:0] n25714_o;
  wire [181:0] n25720_o;
  wire [3:0] n25729_o;
  wire n25739_o;
  wire n25740_o;
  reg [3:0] n25744_q;
  reg [3:0] n25745_q;
  wire n25746_o;
  wire n25747_o;
  wire n25748_o;
  wire n25749_o;
  wire n25752_o;
  wire n25753_o;
  wire n25754_o;
  wire n25755_o;
  reg [150:0] n25758_q;
  reg n25759_q;
  reg n25760_q;
  reg [181:0] n25761_q;
  reg [134:0] n25762_q;
  reg n25763_q;
  reg [2:0] n25764_q;
  reg n25765_q;
  reg [196:0] n25766_q;
  wire n25767_o;
  wire n25768_o;
  reg n25769_q;
  wire [520:0] n25770_o;
  reg [3:0] n25771_q;
  reg n25772_q;
  wire [4:0] n25773_o;
  reg [58:0] n25774_q;
  wire [1:0] n25783_o;
  reg [1:0] n25784_q;
  wire [1:0] n25785_o;
  reg n25787_q;
  reg [47:0] n25788_q;
  reg [1:0] n25789_q;
  wire [67:0] n25790_o;
  wire [66:0] n25791_o;
  localparam [19:0] n25792_o = 20'bZ;
  reg [101:0] n25794_data; // mem_rd
  reg [127:0] n25796_data; // mem_rd
  reg [47:0] n25799_data; // mem_rd
  reg [47:0] n25801_data; // mem_rd
  wire [1:0] n25803_o;
  wire [1:0] n25804_o;
  wire [1:0] n25805_o;
  wire [63:0] n25806_o;
  wire [63:0] n25807_o;
  wire [63:0] n25808_o;
  wire [1:0] n25809_o;
  wire n25810_o;
  wire n25811_o;
  wire n25812_o;
  wire n25813_o;
  wire n25814_o;
  wire n25815_o;
  wire n25816_o;
  wire n25817_o;
  wire n25818_o;
  wire n25819_o;
  wire n25820_o;
  wire n25821_o;
  wire n25822_o;
  wire n25823_o;
  wire n25824_o;
  wire n25825_o;
  wire [3:0] n25826_o;
  wire n25827_o;
  wire n25828_o;
  wire n25829_o;
  wire n25830_o;
  wire n25831_o;
  wire [50:0] n25832_o;
  wire [50:0] n25833_o;
  wire [50:0] n25834_o;
  wire [50:0] n25835_o;
  wire [101:0] n25836_o;
  wire n25837_o;
  wire n25838_o;
  wire [63:0] n25839_o;
  wire [63:0] n25840_o;
  wire [63:0] n25841_o;
  wire [63:0] n25842_o;
  wire [127:0] n25843_o;
  wire [1:0] n25844_o;
  wire n25845_o;
  wire n25846_o;
  wire n25847_o;
  wire n25848_o;
  wire n25849_o;
  wire n25850_o;
  wire n25851_o;
  wire n25852_o;
  wire n25853_o;
  wire n25854_o;
  wire n25855_o;
  wire n25856_o;
  wire n25857_o;
  wire n25858_o;
  wire n25859_o;
  wire n25860_o;
  wire [3:0] n25861_o;
  wire n25862_o;
  wire n25863_o;
  wire n25864_o;
  wire n25865_o;
  wire [1:0] n25866_o;
  reg n25867_o;
  wire n25868_o;
  wire n25869_o;
  wire n25870_o;
  wire n25871_o;
  wire [1:0] n25872_o;
  reg n25873_o;
  wire n25874_o;
  wire n25875_o;
  wire n25876_o;
  wire n25877_o;
  wire n25878_o;
  wire n25879_o;
  wire n25880_o;
  wire n25881_o;
  wire n25882_o;
  wire n25883_o;
  wire n25884_o;
  wire n25885_o;
  wire n25886_o;
  wire [1:0] n25887_o;
  reg n25888_o;
  wire n25889_o;
  wire n25890_o;
  wire n25891_o;
  wire n25892_o;
  wire n25893_o;
  wire n25894_o;
  wire n25895_o;
  wire n25896_o;
  wire [1:0] n25897_o;
  reg n25898_o;
  wire [1:0] n25899_o;
  reg n25900_o;
  wire n25901_o;
  wire n25902_o;
  wire n25903_o;
  wire n25904_o;
  wire n25905_o;
  wire n25906_o;
  wire n25907_o;
  wire n25908_o;
  wire n25909_o;
  wire n25910_o;
  wire n25911_o;
  wire n25912_o;
  wire n25913_o;
  wire n25914_o;
  wire n25915_o;
  wire n25916_o;
  wire n25917_o;
  wire n25918_o;
  wire [3:0] n25919_o;
  wire n25920_o;
  wire n25921_o;
  wire n25922_o;
  wire n25923_o;
  wire n25924_o;
  wire n25925_o;
  wire n25926_o;
  wire n25927_o;
  wire n25928_o;
  wire n25929_o;
  wire n25930_o;
  wire n25931_o;
  wire n25932_o;
  wire n25933_o;
  wire n25934_o;
  wire n25935_o;
  wire n25936_o;
  wire n25937_o;
  wire n25938_o;
  wire n25939_o;
  wire n25940_o;
  wire n25941_o;
  wire n25942_o;
  wire n25943_o;
  wire n25944_o;
  wire n25945_o;
  wire n25946_o;
  wire n25947_o;
  wire n25948_o;
  wire n25949_o;
  wire n25950_o;
  wire n25951_o;
  wire n25952_o;
  wire n25953_o;
  wire [7:0] n25954_o;
  wire n25955_o;
  wire n25956_o;
  wire n25957_o;
  wire n25958_o;
  wire n25959_o;
  wire n25960_o;
  wire n25961_o;
  wire n25962_o;
  wire n25963_o;
  wire n25964_o;
  wire n25965_o;
  wire n25966_o;
  wire n25967_o;
  wire n25968_o;
  wire n25969_o;
  wire n25970_o;
  wire [3:0] n25971_o;
  assign d_out_valid = n23727_o;
  assign d_out_data = n23728_o;
  assign d_out_store_done = n23729_o;
  assign d_out_error = n23730_o;
  assign d_out_cache_paradox = n23731_o;
  assign m_out_stall = n23734_o;
  assign m_out_done = n23735_o;
  assign m_out_err = n23736_o;
  assign m_out_data = n23737_o;
  assign stall_out = r0_stall;
  assign wishbone_out_adr = n23741_o;
  assign wishbone_out_dat = n23742_o;
  assign wishbone_out_sel = n23743_o;
  assign wishbone_out_cyc = n23744_o;
  assign wishbone_out_stb = n23745_o;
  assign wishbone_out_we = n23746_o;
  assign events_load_miss = n23749_o;
  assign events_store_miss = n23750_o;
  assign events_dcache_refill = n23751_o;
  assign events_dtlb_miss = n23752_o;
  assign events_dtlb_miss_resolved = n23753_o;
  assign log_out = n25792_o;
  assign n23725_o = {d_in_byte_sel, d_in_data, d_in_addr, d_in_priv_mode, d_in_virt_mode, d_in_atomic_last, d_in_atomic, d_in_reserve, d_in_nc, d_in_dcbz, d_in_load, d_in_hold, d_in_valid};
  assign n23727_o = n25790_o[0];
  /* mmu.vhdl:23:9  */
  assign n23728_o = n25790_o[64:1];
  /* mmu.vhdl:20:9  */
  assign n23729_o = n25790_o[65];
  /* mmu.vhdl:18:9  */
  assign n23730_o = n25790_o[66];
  assign n23731_o = n25790_o[67];
  assign n23732_o = {m_in_pte, m_in_addr, m_in_tlbld, m_in_doall, m_in_tlbie, m_in_valid};
  /* mmu.vhdl:234:9  */
  assign n23734_o = n25791_o[0];
  assign n23735_o = n25791_o[1];
  /* mmu.vhdl:234:9  */
  assign n23736_o = n25791_o[2];
  assign n23737_o = n25791_o[66:3];
  /* mmu.vhdl:234:9  */
  assign n23738_o = {snoop_in_we, snoop_in_stb, snoop_in_cyc, snoop_in_sel, snoop_in_dat, snoop_in_adr};
  assign n23741_o = n24578_o[28:0];
  /* mmu.vhdl:234:9  */
  assign n23742_o = n24578_o[92:29];
  assign n23743_o = n24578_o[100:93];
  /* mmu.vhdl:234:9  */
  assign n23744_o = n24578_o[101];
  assign n23745_o = n24578_o[102];
  /* mmu.vhdl:234:9  */
  assign n23746_o = n24578_o[103];
  assign n23747_o = {wishbone_in_stall, wishbone_in_ack, wishbone_in_dat};
  assign n23749_o = ev[0];
  assign n23750_o = ev[1];
  assign n23751_o = ev[2];
  assign n23752_o = ev[3];
  assign n23753_o = ev[4];
  /* dcache.vhdl:503:22  */
  assign cache_tag_set = n25801_data; // (signal)
  /* dcache.vhdl:126:12  */
  assign cache_valids = n25744_q; // (signal)
  /* dcache.vhdl:151:12  */
  assign dtlb_valids = n25745_q; // (signal)
  /* dcache.vhdl:283:12  */
  assign r0 = n25758_q; // (signal)
  /* dcache.vhdl:284:12  */
  assign r0_full = n25759_q; // (signal)
  /* dcache.vhdl:354:12  */
  assign r1 = n25770_o; // (signal)
  /* dcache.vhdl:356:12  */
  assign ev = n25773_o; // (signal)
  /* dcache.vhdl:365:12  */
  assign reservation = n25774_q; // (signal)
  /* dcache.vhdl:368:12  */
  assign req_index = n24243_o; // (signal)
  /* dcache.vhdl:369:12  */
  assign req_row = n24252_o; // (signal)
  /* dcache.vhdl:372:12  */
  assign req_op = n24548_o; // (signal)
  /* dcache.vhdl:374:12  */
  assign req_same_tag = n24421_o; // (signal)
  /* dcache.vhdl:375:12  */
  assign req_go = n24267_o; // (signal)
  /* dcache.vhdl:377:12  */
  assign early_req_row = n24570_o; // (signal)
  /* dcache.vhdl:379:12  */
  assign cancel_store = n24605_o; // (signal)
  /* dcache.vhdl:380:12  */
  assign set_rsrv = n24608_o; // (signal)
  /* dcache.vhdl:381:12  */
  assign clear_rsrv = n24611_o; // (signal)
  /* dcache.vhdl:383:12  */
  assign r0_valid = n23854_o; // (signal)
  /* dcache.vhdl:384:12  */
  assign r0_stall = n23848_o; // (signal)
  /* dcache.vhdl:387:12  */
  assign use_forward_st = n24442_o; // (signal)
  /* dcache.vhdl:388:12  */
  assign use_forward_rl = n24445_o; // (signal)
  /* dcache.vhdl:389:12  */
  assign use_forward2 = n24454_o; // (signal)
  /* dcache.vhdl:393:12  */
  assign cache_out = rams_n1_dout; // (signal)
  /* dcache.vhdl:394:12  */
  assign ram_wr_data = n24660_o; // (signal)
  /* dcache.vhdl:395:12  */
  assign ram_wr_select = n24669_o; // (signal)
  /* dcache.vhdl:406:12  */
  assign tlb_tag_way = n25794_data; // (signal)
  /* dcache.vhdl:407:12  */
  assign tlb_pte_way = n25796_data; // (signal)
  /* dcache.vhdl:408:12  */
  assign tlb_valid_way = n25784_q; // (signal)
  /* dcache.vhdl:409:12  */
  assign tlb_req_index = n23916_o; // (signal)
  /* dcache.vhdl:410:12  */
  assign tlb_hit = n23949_o; // (signal)
  /* dcache.vhdl:411:12  */
  assign tlb_hit_way = n23945_o; // (signal)
  /* dcache.vhdl:412:12  */
  assign pte = n23967_o; // (signal)
  /* dcache.vhdl:413:12  */
  assign ra = n24006_o; // (signal)
  /* dcache.vhdl:414:12  */
  assign valid_ra = n23971_o; // (signal)
  /* dcache.vhdl:415:12  */
  assign perm_attr = n24008_o; // (signal)
  /* dcache.vhdl:416:12  */
  assign rc_ok = n24490_o; // (signal)
  /* dcache.vhdl:417:12  */
  assign perm_ok = n24502_o; // (signal)
  /* dcache.vhdl:418:12  */
  assign access_ok = n24504_o; // (signal)
  /* dcache.vhdl:419:12  */
  assign tlb_miss = n23976_o; // (signal)
  /* dcache.vhdl:423:12  */
  assign tlb_plru_victim = n25785_o; // (signal)
  /* dcache.vhdl:503:22  */
  assign snoop_tag_set = n25799_data; // (signal)
  /* dcache.vhdl:426:12  */
  assign snoop_valid = n25787_q; // (signal)
  /* dcache.vhdl:427:12  */
  assign snoop_wrtag = n25788_q; // (signal)
  /* dcache.vhdl:428:12  */
  assign snoop_index = n25789_q; // (signal)
  /* dcache.vhdl:559:18  */
  always @*
    stage_0_r = n23843_q; // (isignal)
  initial
    stage_0_r = 151'bX;
  /* dcache.vhdl:564:21  */
  assign n23761_o = n23732_o[0];
  /* dcache.vhdl:566:41  */
  assign n23763_o = n23732_o[1];
  /* dcache.vhdl:566:55  */
  assign n23764_o = n23732_o[3];
  /* dcache.vhdl:566:47  */
  assign n23765_o = n23763_o | n23764_o;
  /* dcache.vhdl:566:31  */
  assign n23766_o = ~n23765_o;
  /* dcache.vhdl:572:36  */
  assign n23772_o = n23732_o[67:4];
  /* dcache.vhdl:573:36  */
  assign n23773_o = n23732_o[131:68];
  /* dcache.vhdl:575:33  */
  assign n23775_o = n23732_o[1];
  /* dcache.vhdl:576:33  */
  assign n23776_o = n23732_o[2];
  /* dcache.vhdl:577:33  */
  assign n23777_o = n23732_o[3];
  assign n23781_o = n23725_o[145:138];
  /* mmu.vhdl:189:18  */
  assign n23782_o = n23725_o[73:0];
  assign n23788_o = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n23781_o, 64'b0000000000000000000000000000000000000000000000000000000000000000, n23782_o};
  assign n23789_o = {1'b0, 1'b0, 1'b0, n23766_o};
  assign n23790_o = {1'b1, 1'b1, n23777_o, n23776_o, n23775_o, 8'b11111111, n23773_o, n23772_o, 1'b1, 1'b0};
  assign n23791_o = n23788_o[0];
  /* dcache.vhdl:564:13  */
  assign n23792_o = n23761_o ? 1'b1 : n23791_o;
  assign n23793_o = n23788_o[1];
  assign n23794_o = stage_0_r[1];
  /* dcache.vhdl:564:13  */
  assign n23795_o = n23761_o ? n23794_o : n23793_o;
  assign n23796_o = n23788_o[5:2];
  /* dcache.vhdl:564:13  */
  assign n23797_o = n23761_o ? n23789_o : n23796_o;
  assign n23798_o = n23788_o[7:6];
  assign n23799_o = stage_0_r[7:6];
  /* dcache.vhdl:564:13  */
  assign n23800_o = n23761_o ? n23799_o : n23798_o;
  assign n23801_o = n23788_o[150:8];
  /* dcache.vhdl:564:13  */
  assign n23802_o = n23761_o ? n23790_o : n23801_o;
  /* dcache.vhdl:591:23  */
  assign n23803_o = r1[0];
  /* dcache.vhdl:591:28  */
  assign n23804_o = ~n23803_o;
  /* dcache.vhdl:591:43  */
  assign n23805_o = n23725_o[1];
  /* dcache.vhdl:591:48  */
  assign n23806_o = ~n23805_o;
  /* dcache.vhdl:591:34  */
  assign n23807_o = n23804_o & n23806_o;
  /* dcache.vhdl:591:66  */
  assign n23808_o = ~r0_full;
  /* dcache.vhdl:591:55  */
  assign n23809_o = n23807_o | n23808_o;
  assign n23810_o = {n23802_o, n23800_o, n23797_o, n23795_o, n23792_o};
  assign n23811_o = {n23802_o, n23800_o, n23797_o, n23795_o, n23792_o};
  /* dcache.vhdl:593:30  */
  assign n23812_o = n23811_o[145:0];
  /* dcache.vhdl:593:34  */
  assign n23813_o = n23812_o[0];
  /* dcache.vhdl:594:22  */
  assign n23814_o = r0[150];
  /* dcache.vhdl:594:30  */
  assign n23815_o = ~n23814_o;
  /* dcache.vhdl:598:37  */
  assign n23816_o = n23725_o[137:74];
  /* dcache.vhdl:599:34  */
  assign n23817_o = r0[145:0];
  /* dcache.vhdl:599:38  */
  assign n23818_o = n23817_o[0];
  assign n23819_o = r0[137:74];
  /* dcache.vhdl:594:13  */
  assign n23820_o = n23815_o ? n23816_o : n23819_o;
  assign n23821_o = r0[150];
  /* dcache.vhdl:594:13  */
  assign n23822_o = n23815_o ? n23818_o : n23821_o;
  assign n23823_o = n23810_o[73:0];
  assign n23824_o = r0[73:0];
  /* dcache.vhdl:591:13  */
  assign n23825_o = n23809_o ? n23823_o : n23824_o;
  assign n23826_o = n23810_o[137:74];
  /* dcache.vhdl:591:13  */
  assign n23827_o = n23809_o ? n23826_o : n23820_o;
  /* mmu.vhdl:176:5  */
  assign n23828_o = n23810_o[149:138];
  /* mmu.vhdl:177:18  */
  assign n23829_o = r0[149:138];
  /* dcache.vhdl:591:13  */
  assign n23830_o = n23809_o ? n23828_o : n23829_o;
  assign n23831_o = n23810_o[150];
  /* dcache.vhdl:591:13  */
  assign n23832_o = n23809_o ? n23831_o : n23822_o;
  /* dcache.vhdl:591:13  */
  assign n23833_o = n23809_o ? n23813_o : r0_full;
  assign n23834_o = {n23832_o, n23830_o, n23827_o, n23825_o};
  /* dcache.vhdl:589:13  */
  assign n23835_o = rst ? r0 : n23834_o;
  /* dcache.vhdl:589:13  */
  assign n23837_o = rst ? 1'b0 : n23833_o;
  assign n23840_o = {n23802_o, n23800_o, n23797_o, n23795_o, n23792_o};
  /* dcache.vhdl:561:9  */
  always @(posedge clk)
    n23843_q <= n23840_o;
  initial
    n23843_q = 151'bX;
  /* dcache.vhdl:608:33  */
  assign n23845_o = r1[0];
  /* dcache.vhdl:608:46  */
  assign n23846_o = n23725_o[1];
  /* dcache.vhdl:608:38  */
  assign n23847_o = n23845_o | n23846_o;
  /* dcache.vhdl:608:25  */
  assign n23848_o = r0_full & n23847_o;
  /* dcache.vhdl:609:36  */
  assign n23849_o = r1[0];
  /* dcache.vhdl:609:29  */
  assign n23850_o = ~n23849_o;
  /* dcache.vhdl:609:25  */
  assign n23851_o = r0_full & n23850_o;
  /* dcache.vhdl:609:54  */
  assign n23852_o = n23725_o[1];
  /* dcache.vhdl:609:45  */
  assign n23853_o = ~n23852_o;
  /* dcache.vhdl:609:41  */
  assign n23854_o = n23851_o & n23853_o;
  /* dcache.vhdl:622:21  */
  assign n23859_o = n23732_o[0];
  /* dcache.vhdl:623:38  */
  assign n23860_o = n23732_o[16];
  /* dcache.vhdl:625:38  */
  assign n23861_o = n23725_o[22];
  /* dcache.vhdl:622:13  */
  assign n23862_o = n23859_o ? n23860_o : n23861_o;
  /* dcache.vhdl:630:25  */
  assign n23864_o = ~r0_stall;
  /* dcache.vhdl:631:46  */
  assign n23866_o = 1'b1 - n23862_o;
  /* dcache.vhdl:643:20  */
  assign maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_acc = n23896_o; // (signal)
  /* dcache.vhdl:644:20  */
  assign maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_acc_en = n23895_o; // (signal)
  /* dcache.vhdl:645:20  */
  assign maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_out = maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_lru; // (signal)
  /* dcache.vhdl:647:13  */
  plru_1 maybe_tlb_plrus_tlb_plrus_n1_tlb_plru (
    .clk(clk),
    .rst(rst),
    .acc(maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_acc),
    .acc_en(maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_acc_en),
    .lru(maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_lru));
  /* dcache.vhdl:662:23  */
  assign n23889_o = r1[143];
  /* dcache.vhdl:662:37  */
  assign n23890_o = {31'b0, n23889_o};  //  uext
  /* dcache.vhdl:662:37  */
  assign n23892_o = n23890_o == 32'b00000000000000000000000000000000;
  /* dcache.vhdl:663:43  */
  assign n23893_o = r1[141];
  /* dcache.vhdl:662:17  */
  assign n23895_o = n23892_o ? n23893_o : 1'b0;
  /* dcache.vhdl:667:66  */
  assign n23896_o = r1[142];
  /* dcache.vhdl:643:20  */
  assign maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_acc = n23909_o; // (signal)
  /* dcache.vhdl:644:20  */
  assign maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_acc_en = n23908_o; // (signal)
  /* dcache.vhdl:645:20  */
  assign maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_out = maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_lru; // (signal)
  /* dcache.vhdl:647:13  */
  plru_1 maybe_tlb_plrus_tlb_plrus_n2_tlb_plru (
    .clk(clk),
    .rst(rst),
    .acc(maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_acc),
    .acc_en(maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_acc_en),
    .lru(maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_lru));
  /* dcache.vhdl:662:23  */
  assign n23902_o = r1[143];
  /* dcache.vhdl:662:37  */
  assign n23903_o = {31'b0, n23902_o};  //  uext
  /* dcache.vhdl:662:37  */
  assign n23905_o = n23903_o == 32'b00000000000000000000000000000001;
  /* dcache.vhdl:663:43  */
  assign n23906_o = r1[141];
  /* dcache.vhdl:662:17  */
  assign n23908_o = n23905_o ? n23906_o : 1'b0;
  /* dcache.vhdl:667:66  */
  assign n23909_o = r1[142];
  /* dcache.vhdl:678:57  */
  assign n23916_o = r0[22];
  /* dcache.vhdl:682:29  */
  assign n23918_o = r0[73:23];
  /* dcache.vhdl:684:29  */
  assign n23919_o = tlb_valid_way[0];
  /* dcache.vhdl:511:20  */
  assign n23926_o = tlb_tag_way[50:0];
  /* dcache.vhdl:685:46  */
  assign n23927_o = n23926_o == n23918_o;
  /* dcache.vhdl:684:39  */
  assign n23928_o = n23919_o & n23927_o;
  /* dcache.vhdl:684:13  */
  assign n23931_o = n23928_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:684:29  */
  assign n23933_o = tlb_valid_way[1];
  /* dcache.vhdl:511:20  */
  assign n23940_o = tlb_tag_way[101:51];
  /* dcache.vhdl:685:46  */
  assign n23941_o = n23940_o == n23918_o;
  /* dcache.vhdl:684:39  */
  assign n23942_o = n23933_o & n23941_o;
  /* dcache.vhdl:684:13  */
  assign n23945_o = n23942_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:684:13  */
  assign n23948_o = n23942_o ? 1'b1 : n23931_o;
  /* dcache.vhdl:690:24  */
  assign n23949_o = n23948_o & r0_valid;
  /* dcache.vhdl:692:9  */
  assign n23967_o = tlb_hit ? n25808_o : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* dcache.vhdl:697:39  */
  assign n23968_o = r0[145:0];
  /* dcache.vhdl:697:43  */
  assign n23969_o = n23968_o[8];
  /* dcache.vhdl:697:32  */
  assign n23970_o = ~n23969_o;
  /* dcache.vhdl:697:29  */
  assign n23971_o = tlb_hit | n23970_o;
  /* dcache.vhdl:698:37  */
  assign n23972_o = r0[145:0];
  /* dcache.vhdl:698:41  */
  assign n23973_o = n23972_o[8];
  /* dcache.vhdl:698:30  */
  assign n23974_o = r0_valid & n23973_o;
  /* dcache.vhdl:698:55  */
  assign n23975_o = ~tlb_hit;
  /* dcache.vhdl:698:51  */
  assign n23976_o = n23974_o & n23975_o;
  /* dcache.vhdl:699:15  */
  assign n23977_o = r0[145:0];
  /* dcache.vhdl:699:19  */
  assign n23978_o = n23977_o[8];
  /* dcache.vhdl:700:22  */
  assign n23979_o = pte[55:12];
  /* dcache.vhdl:701:30  */
  assign n23980_o = r0[21:13];
  /* dcache.vhdl:700:62  */
  assign n23981_o = {n23979_o, n23980_o};
  /* dcache.vhdl:701:68  */
  assign n23983_o = {n23981_o, 3'b000};
  /* dcache.vhdl:170:28  */
  assign n23990_o = pte[8];
  /* dcache.vhdl:171:26  */
  assign n23993_o = pte[7];
  /* dcache.vhdl:172:26  */
  assign n23995_o = pte[5];
  /* dcache.vhdl:173:23  */
  assign n23997_o = pte[3];
  /* dcache.vhdl:174:26  */
  assign n23999_o = pte[2];
  /* dcache.vhdl:175:26  */
  assign n24001_o = pte[1];
  assign n24002_o = {n24001_o, n23999_o, n23997_o, n23995_o, n23993_o, n23990_o};
  /* dcache.vhdl:705:30  */
  assign n24003_o = r0[65:13];
  /* dcache.vhdl:705:71  */
  assign n24005_o = {n24003_o, 3'b000};
  /* dcache.vhdl:699:9  */
  assign n24006_o = n23978_o ? n23983_o : n24005_o;
  /* dcache.vhdl:699:9  */
  assign n24008_o = n23978_o ? n24002_o : 6'b111011;
  /* dcache.vhdl:720:38  */
  assign n24019_o = r0[146];
  /* dcache.vhdl:720:31  */
  assign n24020_o = r0_valid & n24019_o;
  /* dcache.vhdl:721:38  */
  assign n24021_o = r0[148];
  /* dcache.vhdl:721:31  */
  assign n24022_o = r0_valid & n24021_o;
  /* dcache.vhdl:723:49  */
  assign n24023_o = r0[147];
  /* dcache.vhdl:723:42  */
  assign n24024_o = n24020_o & n24023_o;
  /* dcache.vhdl:723:26  */
  assign n24025_o = rst | n24024_o;
  /* dcache.vhdl:730:33  */
  assign n24029_o = 1'b1 - tlb_req_index;
  /* dcache.vhdl:729:17  */
  assign n24035_o = tlb_hit ? n25826_o : dtlb_valids;
  /* dcache.vhdl:736:69  */
  assign n24037_o = 1'b1 - tlb_req_index;
  /* dcache.vhdl:733:17  */
  assign n24041_o = tlb_hit ? tlb_hit_way : n25829_o;
  /* dcache.vhdl:738:37  */
  assign n24042_o = r0[73:23];
  /* dcache.vhdl:743:52  */
  assign n24062_o = r0[145:0];
  /* dcache.vhdl:743:56  */
  assign n24063_o = n24062_o[137:74];
  /* dcache.vhdl:745:29  */
  assign n24082_o = 1'b1 - tlb_req_index;
  /* dcache.vhdl:732:13  */
  assign n24088_o = n24022_o ? n25861_o : dtlb_valids;
  /* dcache.vhdl:728:13  */
  assign n24095_o = n24020_o ? n24035_o : n24088_o;
  assign n24102_o = {2'b00, 2'b00};
  /* dcache.vhdl:723:13  */
  assign n24103_o = n24025_o ? n24102_o : n24095_o;
  /* dcache.vhdl:793:24  */
  assign n24129_o = n23732_o[0];
  /* dcache.vhdl:794:41  */
  assign n24131_o = n23732_o[67:4];
  /* dcache.vhdl:437:40  */
  assign n24136_o = n24131_o[7:6];
  /* dcache.vhdl:796:41  */
  assign n24139_o = n23725_o[73:10];
  /* dcache.vhdl:437:40  */
  assign n24144_o = n24139_o[7:6];
  /* dcache.vhdl:793:13  */
  assign n24146_o = n24129_o ? n24136_o : n24144_o;
  /* dcache.vhdl:791:13  */
  assign n24147_o = r0_stall ? req_index : n24146_o;
  /* dcache.vhdl:807:54  */
  assign n24160_o = n23738_o[28:0];
  assign n24167_o = n24166_o[63:32];
  assign n24168_o = n24166_o[2:0];
  assign n24169_o = {n24167_o, n24160_o, n24168_o};
  /* common.vhdl:790:20  */
  assign n24174_o = n24169_o[55:0];
  /* dcache.vhdl:437:40  */
  assign n24180_o = n24174_o[7:6];
  /* dcache.vhdl:497:20  */
  assign n24191_o = n24174_o[55:8];
  /* dcache.vhdl:437:40  */
  assign n24197_o = n24174_o[7:6];
  /* dcache.vhdl:813:24  */
  assign n24199_o = r1[443:340];
  /* dcache.vhdl:813:27  */
  assign n24200_o = n24199_o[101];
  /* dcache.vhdl:813:53  */
  assign n24201_o = n23747_o[65];
  /* dcache.vhdl:813:59  */
  assign n24202_o = ~n24201_o;
  /* dcache.vhdl:813:37  */
  assign n24203_o = n24200_o & n24202_o;
  /* dcache.vhdl:813:16  */
  assign n24204_o = ~n24203_o;
  /* dcache.vhdl:814:41  */
  assign n24205_o = n23738_o[101];
  /* dcache.vhdl:814:58  */
  assign n24206_o = n23738_o[102];
  /* dcache.vhdl:814:45  */
  assign n24207_o = n24205_o & n24206_o;
  /* dcache.vhdl:814:75  */
  assign n24208_o = n23738_o[103];
  /* dcache.vhdl:814:62  */
  assign n24209_o = n24207_o & n24208_o;
  /* dcache.vhdl:813:13  */
  assign n24211_o = n24204_o ? n24209_o : 1'b0;
  /* dcache.vhdl:839:35  */
  assign n24237_o = r0[145:0];
  /* dcache.vhdl:839:39  */
  assign n24238_o = n24237_o[73:10];
  /* dcache.vhdl:437:40  */
  assign n24243_o = n24238_o[7:6];
  /* dcache.vhdl:840:31  */
  assign n24246_o = r0[145:0];
  /* dcache.vhdl:840:35  */
  assign n24247_o = n24246_o[73:10];
  /* dcache.vhdl:443:40  */
  assign n24252_o = n24247_o[7:3];
  /* dcache.vhdl:843:36  */
  assign n24260_o = r0[146];
  /* dcache.vhdl:843:48  */
  assign n24261_o = r0[148];
  /* dcache.vhdl:843:42  */
  assign n24262_o = n24260_o | n24261_o;
  /* dcache.vhdl:843:28  */
  assign n24263_o = ~n24262_o;
  /* dcache.vhdl:843:24  */
  assign n24264_o = r0_valid & n24263_o;
  /* dcache.vhdl:843:66  */
  assign n24265_o = r1[516];
  /* dcache.vhdl:843:59  */
  assign n24266_o = ~n24265_o;
  /* dcache.vhdl:843:55  */
  assign n24267_o = n24264_o & n24266_o;
  /* dcache.vhdl:853:15  */
  assign n24268_o = r0[145:0];
  /* dcache.vhdl:853:19  */
  assign n24269_o = n24268_o[8];
  /* dcache.vhdl:528:20  */
  assign n24276_o = tlb_pte_way[63:0];
  /* dcache.vhdl:860:30  */
  assign n24277_o = n24276_o[55:12];
  /* dcache.vhdl:861:36  */
  assign n24278_o = r0[21:10];
  /* dcache.vhdl:860:70  */
  assign n24279_o = {n24277_o, n24278_o};
  /* dcache.vhdl:497:20  */
  assign n24285_o = n24279_o[55:8];
  /* dcache.vhdl:864:50  */
  assign n24287_o = 2'b11 - req_index;
  /* dcache.vhdl:864:33  */
  assign n24290_o = n24267_o & n25867_o;
  /* dcache.vhdl:865:52  */
  assign n24296_o = cache_tag_set == n24285_o;
  /* dcache.vhdl:864:70  */
  assign n24297_o = n24290_o & n24296_o;
  /* dcache.vhdl:866:38  */
  assign n24298_o = tlb_valid_way[0];
  /* dcache.vhdl:865:60  */
  assign n24299_o = n24297_o & n24298_o;
  /* dcache.vhdl:864:21  */
  assign n24302_o = n24299_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:872:31  */
  assign n24304_o = r1[491:444];
  /* dcache.vhdl:872:26  */
  assign n24305_o = n24285_o == n24304_o;
  /* dcache.vhdl:872:17  */
  assign n24308_o = n24305_o ? 1'b1 : 1'b0;
  assign n24310_o = n24309_o[1];
  /* dcache.vhdl:875:31  */
  assign n24311_o = r1[255:208];
  /* dcache.vhdl:875:26  */
  assign n24312_o = n24285_o == n24311_o;
  /* dcache.vhdl:875:17  */
  assign n24315_o = n24312_o ? 1'b1 : 1'b0;
  assign n24317_o = n24316_o[1];
  /* dcache.vhdl:528:20  */
  assign n24324_o = tlb_pte_way[127:64];
  /* dcache.vhdl:860:30  */
  assign n24325_o = n24324_o[55:12];
  /* dcache.vhdl:861:36  */
  assign n24326_o = r0[21:10];
  /* dcache.vhdl:860:70  */
  assign n24327_o = {n24325_o, n24326_o};
  /* dcache.vhdl:497:20  */
  assign n24333_o = n24327_o[55:8];
  /* dcache.vhdl:864:50  */
  assign n24335_o = 2'b11 - req_index;
  /* dcache.vhdl:864:33  */
  assign n24338_o = n24267_o & n25873_o;
  /* dcache.vhdl:865:52  */
  assign n24344_o = cache_tag_set == n24333_o;
  /* dcache.vhdl:864:70  */
  assign n24345_o = n24338_o & n24344_o;
  /* dcache.vhdl:866:38  */
  assign n24346_o = tlb_valid_way[1];
  /* dcache.vhdl:865:60  */
  assign n24347_o = n24345_o & n24346_o;
  /* dcache.vhdl:864:21  */
  assign n24350_o = n24347_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:872:31  */
  assign n24352_o = r1[491:444];
  /* dcache.vhdl:872:26  */
  assign n24353_o = n24333_o == n24352_o;
  /* dcache.vhdl:872:17  */
  assign n24355_o = n24353_o ? 1'b1 : n24310_o;
  /* dcache.vhdl:875:31  */
  assign n24356_o = r1[255:208];
  /* dcache.vhdl:875:26  */
  assign n24357_o = n24333_o == n24356_o;
  /* dcache.vhdl:875:17  */
  assign n24359_o = n24357_o ? 1'b1 : n24317_o;
  /* dcache.vhdl:880:34  */
  assign n24361_o = {n24350_o, n24302_o};
  /* dcache.vhdl:882:41  */
  assign n24367_o = {n24355_o, n24308_o};
  /* dcache.vhdl:883:41  */
  assign n24370_o = {n24359_o, n24315_o};
  /* dcache.vhdl:879:13  */
  assign n24373_o = tlb_hit ? n25876_o : 1'b0;
  /* dcache.vhdl:879:13  */
  assign n24375_o = tlb_hit ? n25879_o : 1'b0;
  /* dcache.vhdl:879:13  */
  assign n24377_o = tlb_hit ? n25882_o : 1'b0;
  /* dcache.vhdl:886:33  */
  assign n24379_o = r0[145:0];
  /* dcache.vhdl:886:37  */
  assign n24380_o = n24379_o[73:10];
  /* dcache.vhdl:497:20  */
  assign n24385_o = n24380_o[55:8];
  /* dcache.vhdl:888:46  */
  assign n24387_o = 2'b11 - req_index;
  /* dcache.vhdl:888:29  */
  assign n24390_o = n24267_o & n25888_o;
  /* dcache.vhdl:889:48  */
  assign n24396_o = cache_tag_set == n24385_o;
  /* dcache.vhdl:888:66  */
  assign n24397_o = n24390_o & n24396_o;
  /* dcache.vhdl:888:17  */
  assign n24400_o = n24397_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:894:27  */
  assign n24401_o = r1[491:444];
  /* dcache.vhdl:894:22  */
  assign n24402_o = n24385_o == n24401_o;
  /* dcache.vhdl:894:13  */
  assign n24405_o = n24402_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:897:27  */
  assign n24406_o = r1[255:208];
  /* dcache.vhdl:897:22  */
  assign n24407_o = n24385_o == n24406_o;
  /* dcache.vhdl:897:13  */
  assign n24410_o = n24407_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:853:9  */
  assign n24411_o = n24269_o ? n24373_o : n24400_o;
  /* dcache.vhdl:853:9  */
  assign n24421_o = n24269_o ? n24375_o : n24405_o;
  /* dcache.vhdl:853:9  */
  assign n24425_o = n24269_o ? n24377_o : n24410_o;
  /* dcache.vhdl:907:15  */
  assign n24427_o = r1[496:492];
  /* dcache.vhdl:907:25  */
  assign n24428_o = {27'b0, n24427_o};  //  uext
  /* dcache.vhdl:907:25  */
  assign n24429_o = {27'b0, req_row};  //  uext
  /* dcache.vhdl:907:25  */
  assign n24430_o = n24428_o == n24429_o;
  /* dcache.vhdl:907:35  */
  assign n24431_o = n24430_o & n24421_o;
  /* dcache.vhdl:909:34  */
  assign n24432_o = r1[337];
  /* dcache.vhdl:910:19  */
  assign n24433_o = r1[335:334];
  /* dcache.vhdl:910:25  */
  assign n24435_o = n24433_o == 2'b01;
  /* dcache.vhdl:910:59  */
  assign n24436_o = n23747_o[64];
  /* dcache.vhdl:910:43  */
  assign n24437_o = n24435_o & n24436_o;
  /* dcache.vhdl:910:13  */
  assign n24440_o = n24437_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:907:9  */
  assign n24442_o = n24431_o ? n24432_o : 1'b0;
  /* dcache.vhdl:907:9  */
  assign n24445_o = n24431_o ? n24440_o : 1'b0;
  /* dcache.vhdl:915:15  */
  assign n24447_o = r1[269:265];
  /* dcache.vhdl:915:27  */
  assign n24448_o = {27'b0, n24447_o};  //  uext
  /* dcache.vhdl:915:27  */
  assign n24449_o = {27'b0, req_row};  //  uext
  /* dcache.vhdl:915:27  */
  assign n24450_o = n24448_o == n24449_o;
  /* dcache.vhdl:915:37  */
  assign n24451_o = n24450_o & n24425_o;
  /* dcache.vhdl:916:32  */
  assign n24452_o = r1[264];
  /* dcache.vhdl:915:9  */
  assign n24454_o = n24451_o ? n24452_o : 1'b0;
  /* dcache.vhdl:927:15  */
  assign n24463_o = r1[335:334];
  /* dcache.vhdl:927:21  */
  assign n24465_o = n24463_o == 2'b01;
  /* dcache.vhdl:927:53  */
  assign n24466_o = {30'b0, req_index};  //  uext
  /* dcache.vhdl:927:58  */
  assign n24467_o = r1[498:497];
  /* dcache.vhdl:927:53  */
  assign n24468_o = {30'b0, n24467_o};  //  uext
  /* dcache.vhdl:927:53  */
  assign n24469_o = n24466_o == n24468_o;
  /* dcache.vhdl:927:39  */
  assign n24470_o = n24465_o & n24469_o;
  /* dcache.vhdl:927:70  */
  assign n24471_o = n24470_o & n24421_o;
  /* dcache.vhdl:935:30  */
  assign n24472_o = r0[145:0];
  /* dcache.vhdl:935:34  */
  assign n24473_o = n24472_o[2];
  /* dcache.vhdl:935:23  */
  assign n24474_o = ~n24473_o;
  /* dcache.vhdl:935:64  */
  assign n24475_o = {27'b0, req_row};  //  uext
  assign n24476_o = n24475_o[2:0];
  /* dcache.vhdl:935:64  */
  assign n24479_o = 3'b111 - n24476_o;
  /* dcache.vhdl:935:39  */
  assign n24482_o = n24474_o | n25902_o;
  /* dcache.vhdl:935:82  */
  assign n24483_o = n24482_o | use_forward_rl;
  /* dcache.vhdl:927:9  */
  assign n24484_o = n24471_o ? n24483_o : n24411_o;
  /* dcache.vhdl:945:28  */
  assign n24485_o = perm_attr[0];
  /* dcache.vhdl:945:46  */
  assign n24486_o = r0[145:0];
  /* dcache.vhdl:945:50  */
  assign n24487_o = n24486_o[2];
  /* dcache.vhdl:945:68  */
  assign n24488_o = perm_attr[1];
  /* dcache.vhdl:945:55  */
  assign n24489_o = n24487_o | n24488_o;
  /* dcache.vhdl:945:38  */
  assign n24490_o = n24485_o & n24489_o;
  /* dcache.vhdl:946:24  */
  assign n24491_o = r0[145:0];
  /* dcache.vhdl:946:28  */
  assign n24492_o = n24491_o[9];
  /* dcache.vhdl:946:55  */
  assign n24493_o = perm_attr[3];
  /* dcache.vhdl:946:41  */
  assign n24494_o = ~n24493_o;
  /* dcache.vhdl:946:38  */
  assign n24495_o = n24492_o | n24494_o;
  /* dcache.vhdl:947:31  */
  assign n24496_o = perm_attr[5];
  /* dcache.vhdl:947:46  */
  assign n24497_o = r0[145:0];
  /* dcache.vhdl:947:50  */
  assign n24498_o = n24497_o[2];
  /* dcache.vhdl:947:69  */
  assign n24499_o = perm_attr[4];
  /* dcache.vhdl:947:55  */
  assign n24500_o = n24498_o & n24499_o;
  /* dcache.vhdl:947:39  */
  assign n24501_o = n24496_o | n24500_o;
  /* dcache.vhdl:946:61  */
  assign n24502_o = n24495_o & n24501_o;
  /* dcache.vhdl:948:31  */
  assign n24503_o = valid_ra & perm_ok;
  /* dcache.vhdl:948:43  */
  assign n24504_o = n24503_o & rc_ok;
  /* dcache.vhdl:953:18  */
  assign n24505_o = r0[145:0];
  /* dcache.vhdl:953:22  */
  assign n24506_o = n24505_o[4];
  /* dcache.vhdl:953:38  */
  assign n24507_o = perm_attr[2];
  /* dcache.vhdl:953:25  */
  assign n24508_o = n24506_o | n24507_o;
  /* dcache.vhdl:956:26  */
  assign n24509_o = ~access_ok;
  /* dcache.vhdl:961:29  */
  assign n24510_o = r0[145:0];
  /* dcache.vhdl:961:33  */
  assign n24511_o = n24510_o[2];
  /* dcache.vhdl:961:38  */
  assign n24512_o = {n24511_o, n24508_o};
  /* dcache.vhdl:961:43  */
  assign n24513_o = {n24512_o, n24484_o};
  /* dcache.vhdl:963:21  */
  assign n24515_o = n24513_o == 3'b101;
  /* dcache.vhdl:964:21  */
  assign n24517_o = n24513_o == 3'b100;
  /* dcache.vhdl:965:21  */
  assign n24519_o = n24513_o == 3'b110;
  /* dcache.vhdl:966:21  */
  assign n24521_o = n24513_o == 3'b001;
  /* dcache.vhdl:967:21  */
  assign n24523_o = n24513_o == 3'b000;
  /* dcache.vhdl:968:21  */
  assign n24525_o = n24513_o == 3'b010;
  /* dcache.vhdl:969:21  */
  assign n24527_o = n24513_o == 3'b011;
  /* dcache.vhdl:970:21  */
  assign n24529_o = n24513_o == 3'b111;
  assign n24530_o = {n24529_o, n24527_o, n24525_o, n24523_o, n24521_o, n24519_o, n24517_o, n24515_o};
  /* dcache.vhdl:962:17  */
  always @*
    case (n24530_o)
      8'b10000000: n24540_o = 3'b001;
      8'b01000000: n24540_o = 3'b001;
      8'b00100000: n24540_o = 3'b111;
      8'b00010000: n24540_o = 3'b111;
      8'b00001000: n24540_o = 3'b110;
      8'b00000100: n24540_o = 3'b101;
      8'b00000010: n24540_o = 3'b100;
      8'b00000001: n24540_o = 3'b011;
      default: n24540_o = 3'b000;
    endcase
  /* dcache.vhdl:958:13  */
  assign n24542_o = cancel_store ? 3'b010 : n24540_o;
  /* dcache.vhdl:956:13  */
  assign n24545_o = n24509_o ? 3'b001 : n24542_o;
  /* dcache.vhdl:955:9  */
  assign n24548_o = n24267_o ? n24545_o : 3'b000;
  /* dcache.vhdl:982:21  */
  assign n24551_o = ~r0_stall;
  /* dcache.vhdl:983:21  */
  assign n24552_o = n23732_o[0];
  /* dcache.vhdl:984:47  */
  assign n24554_o = n23732_o[67:4];
  /* dcache.vhdl:443:40  */
  assign n24559_o = n24554_o[7:3];
  /* dcache.vhdl:986:47  */
  assign n24562_o = n23725_o[73:10];
  /* dcache.vhdl:443:40  */
  assign n24567_o = n24562_o[7:3];
  /* dcache.vhdl:983:13  */
  assign n24569_o = n24552_o ? n24559_o : n24567_o;
  /* dcache.vhdl:982:9  */
  assign n24570_o = n24551_o ? n24569_o : req_row;
  /* dcache.vhdl:994:24  */
  assign n24578_o = r1[443:340];
  /* dcache.vhdl:1002:34  */
  assign n24580_o = r0[145:0];
  /* dcache.vhdl:1002:38  */
  assign n24581_o = n24580_o[5];
  /* dcache.vhdl:1002:27  */
  assign n24582_o = r0_valid & n24581_o;
  /* dcache.vhdl:1005:19  */
  assign n24583_o = r0[145:0];
  /* dcache.vhdl:1005:23  */
  assign n24584_o = n24583_o[2];
  /* dcache.vhdl:1007:32  */
  assign n24585_o = r0[145:0];
  /* dcache.vhdl:1007:36  */
  assign n24586_o = n24585_o[7];
  /* dcache.vhdl:1010:34  */
  assign n24587_o = r0[145:0];
  /* dcache.vhdl:1010:38  */
  assign n24588_o = n24587_o[7];
  /* dcache.vhdl:1011:32  */
  assign n24589_o = reservation[0];
  /* dcache.vhdl:1011:38  */
  assign n24590_o = ~n24589_o;
  /* dcache.vhdl:1012:32  */
  assign n24591_o = r0[73:16];
  /* dcache.vhdl:1012:73  */
  assign n24592_o = reservation[58:1];
  /* dcache.vhdl:1012:58  */
  assign n24593_o = n24591_o != n24592_o;
  /* dcache.vhdl:1011:44  */
  assign n24594_o = n24590_o | n24593_o;
  /* dcache.vhdl:1011:17  */
  assign n24597_o = n24594_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:1005:13  */
  assign n24599_o = n24584_o ? 1'b0 : n24597_o;
  /* dcache.vhdl:1005:13  */
  assign n24601_o = n24584_o ? n24586_o : 1'b0;
  /* dcache.vhdl:1005:13  */
  assign n24603_o = n24584_o ? 1'b0 : n24588_o;
  /* dcache.vhdl:1002:9  */
  assign n24605_o = n24582_o ? n24599_o : 1'b0;
  /* dcache.vhdl:1002:9  */
  assign n24608_o = n24582_o ? n24601_o : 1'b0;
  /* dcache.vhdl:1002:9  */
  assign n24611_o = n24582_o ? n24603_o : 1'b0;
  /* dcache.vhdl:1024:34  */
  assign n24617_o = r0_valid & access_ok;
  /* dcache.vhdl:1029:52  */
  assign n24620_o = r0[73:16];
  assign n24621_o = {n24620_o, 1'b1};
  /* dcache.vhdl:1027:17  */
  assign n24622_o = set_rsrv ? n24621_o : reservation;
  assign n24623_o = n24622_o[0];
  /* dcache.vhdl:1025:17  */
  assign n24624_o = clear_rsrv ? 1'b0 : n24623_o;
  assign n24625_o = n24622_o[58:1];
  assign n24626_o = reservation[58:1];
  /* dcache.vhdl:1025:17  */
  assign n24627_o = clear_rsrv ? n24626_o : n24625_o;
  assign n24628_o = {n24627_o, n24624_o};
  /* dcache.vhdl:1024:13  */
  assign n24629_o = n24617_o ? n24628_o : reservation;
  assign n24630_o = n24629_o[0];
  /* dcache.vhdl:1022:13  */
  assign n24631_o = rst ? 1'b0 : n24630_o;
  assign n24632_o = n24629_o[58:1];
  assign n24633_o = reservation[58:1];
  /* dcache.vhdl:1022:13  */
  assign n24634_o = rst ? n24633_o : n24632_o;
  assign n24635_o = {n24634_o, n24631_o};
  /* dcache.vhdl:1039:27  */
  assign n24639_o = r1[515];
  /* dcache.vhdl:1040:26  */
  assign n24640_o = r1[333:270];
  /* dcache.vhdl:1041:36  */
  assign n24641_o = r1[520];
  /* dcache.vhdl:1041:29  */
  assign n24642_o = ~n24641_o;
  /* dcache.vhdl:1042:27  */
  assign n24643_o = r1[516];
  /* dcache.vhdl:1043:35  */
  assign n24644_o = r1[519];
  /* dcache.vhdl:1046:26  */
  assign n24645_o = r1[517];
  /* dcache.vhdl:1047:25  */
  assign n24646_o = r1[518];
  /* dcache.vhdl:1048:26  */
  assign n24647_o = r1[333:270];
  /* dcache.vhdl:1105:23  */
  assign n24657_o = r1[136:2];
  /* dcache.vhdl:1105:27  */
  assign n24658_o = n24657_o[124:61];
  /* dcache.vhdl:1105:40  */
  assign n24659_o = r1[337];
  /* dcache.vhdl:1105:32  */
  assign n24660_o = n24659_o ? n24658_o : n24664_o;
  /* dcache.vhdl:1106:32  */
  assign n24661_o = n23747_o[63:0];
  /* dcache.vhdl:1106:44  */
  assign n24662_o = r1[336];
  /* dcache.vhdl:1106:49  */
  assign n24663_o = ~n24662_o;
  /* dcache.vhdl:1105:57  */
  assign n24664_o = n24663_o ? n24661_o : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* dcache.vhdl:1108:25  */
  assign n24666_o = r1[136:2];
  /* dcache.vhdl:1108:29  */
  assign n24667_o = n24666_o[132:125];
  /* dcache.vhdl:1108:46  */
  assign n24668_o = r1[337];
  /* dcache.vhdl:1108:38  */
  assign n24669_o = n24668_o ? n24667_o : 8'b11111111;
  /* dcache.vhdl:1122:16  */
  assign rams_n1_do_read = 1'b1; // (signal)
  /* dcache.vhdl:1123:16  */
  assign rams_n1_rd_addr = early_req_row; // (signal)
  /* dcache.vhdl:1125:16  */
  assign rams_n1_wr_addr = n24675_o; // (signal)
  /* dcache.vhdl:1128:16  */
  assign rams_n1_wr_sel_m = n24687_o; // (signal)
  /* dcache.vhdl:1129:16  */
  assign rams_n1_dout = rams_n1_way_rd_data; // (signal)
  /* dcache.vhdl:1131:9  */
  cache_ram_5_64_1489f923c4dca729178b3e3233458550d8dddf29 rams_n1_way (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(clk),
    .rd_en(rams_n1_do_read),
    .rd_addr(rams_n1_rd_addr),
    .wr_sel(rams_n1_wr_sel_m),
    .wr_addr(rams_n1_wr_addr),
    .wr_data(ram_wr_data),
    .rd_data(rams_n1_way_rd_data));
  /* dcache.vhdl:1160:57  */
  assign n24675_o = r1[496:492];
  /* dcache.vhdl:1164:21  */
  assign n24677_o = r1[337];
  /* dcache.vhdl:1165:22  */
  assign n24678_o = r1[335:334];
  /* dcache.vhdl:1165:28  */
  assign n24680_o = n24678_o == 2'b01;
  /* dcache.vhdl:1165:62  */
  assign n24681_o = n23747_o[64];
  /* dcache.vhdl:1165:46  */
  assign n24682_o = n24680_o & n24681_o;
  /* dcache.vhdl:1164:38  */
  assign n24683_o = n24677_o | n24682_o;
  /* dcache.vhdl:1163:32  */
  assign n24685_o = 1'b1 & n24683_o;
  /* dcache.vhdl:1163:13  */
  assign n24687_o = n24685_o ? ram_wr_select : 8'b00000000;
  /* dcache.vhdl:1191:34  */
  assign n24701_o = r0[149];
  /* dcache.vhdl:1199:23  */
  assign n24704_o = r1[0];
  /* dcache.vhdl:1199:34  */
  assign n24705_o = n24704_o | use_forward_rl;
  /* dcache.vhdl:1200:37  */
  assign n24706_o = r1[336];
  /* dcache.vhdl:1200:32  */
  assign n24708_o = {1'b0, n24706_o};
  /* dcache.vhdl:1201:63  */
  assign n24709_o = r1[127];
  /* dcache.vhdl:1201:44  */
  assign n24710_o = use_forward_st & n24709_o;
  /* dcache.vhdl:1203:60  */
  assign n24711_o = r1[256];
  /* dcache.vhdl:1203:42  */
  assign n24712_o = use_forward2 & n24711_o;
  /* dcache.vhdl:1203:17  */
  assign n24715_o = n24712_o ? 2'b10 : 2'b11;
  /* dcache.vhdl:1201:17  */
  assign n24717_o = n24710_o ? 2'b01 : n24715_o;
  /* dcache.vhdl:1199:17  */
  assign n24718_o = n24705_o ? n24708_o : n24717_o;
  /* dcache.vhdl:1211:68  */
  assign n24719_o = n23747_o[7:0];
  /* dcache.vhdl:1210:21  */
  assign n24721_o = n24718_o == 2'b00;
  /* dcache.vhdl:1213:64  */
  assign n24722_o = r1[70:63];
  /* dcache.vhdl:1212:21  */
  assign n24724_o = n24718_o == 2'b01;
  /* dcache.vhdl:1215:68  */
  assign n24725_o = r1[151:144];
  /* dcache.vhdl:1214:21  */
  assign n24727_o = n24718_o == 2'b10;
  /* dcache.vhdl:1217:75  */
  assign n24728_o = cache_out[7:0];
  assign n24729_o = {n24727_o, n24724_o, n24721_o};
  /* dcache.vhdl:1209:17  */
  always @*
    case (n24729_o)
      3'b100: n24730_o = n24725_o;
      3'b010: n24730_o = n24722_o;
      3'b001: n24730_o = n24719_o;
      default: n24730_o = n24728_o;
    endcase
  /* dcache.vhdl:1199:23  */
  assign n24731_o = r1[0];
  /* dcache.vhdl:1199:34  */
  assign n24732_o = n24731_o | use_forward_rl;
  /* dcache.vhdl:1200:37  */
  assign n24733_o = r1[336];
  /* dcache.vhdl:1200:32  */
  assign n24735_o = {1'b0, n24733_o};
  /* dcache.vhdl:1201:63  */
  assign n24736_o = r1[128];
  /* dcache.vhdl:1201:44  */
  assign n24737_o = use_forward_st & n24736_o;
  /* dcache.vhdl:1203:60  */
  assign n24738_o = r1[257];
  /* dcache.vhdl:1203:42  */
  assign n24739_o = use_forward2 & n24738_o;
  /* dcache.vhdl:1203:17  */
  assign n24742_o = n24739_o ? 2'b10 : 2'b11;
  /* dcache.vhdl:1201:17  */
  assign n24744_o = n24737_o ? 2'b01 : n24742_o;
  /* dcache.vhdl:1199:17  */
  assign n24745_o = n24732_o ? n24735_o : n24744_o;
  /* dcache.vhdl:1211:68  */
  assign n24746_o = n23747_o[15:8];
  /* dcache.vhdl:1210:21  */
  assign n24748_o = n24745_o == 2'b00;
  /* dcache.vhdl:1213:64  */
  assign n24749_o = r1[78:71];
  /* dcache.vhdl:1212:21  */
  assign n24751_o = n24745_o == 2'b01;
  /* dcache.vhdl:1215:68  */
  assign n24752_o = r1[159:152];
  /* dcache.vhdl:1214:21  */
  assign n24754_o = n24745_o == 2'b10;
  /* dcache.vhdl:1217:75  */
  assign n24755_o = cache_out[15:8];
  assign n24756_o = {n24754_o, n24751_o, n24748_o};
  /* dcache.vhdl:1209:17  */
  always @*
    case (n24756_o)
      3'b100: n24757_o = n24752_o;
      3'b010: n24757_o = n24749_o;
      3'b001: n24757_o = n24746_o;
      default: n24757_o = n24755_o;
    endcase
  /* dcache.vhdl:1199:23  */
  assign n24758_o = r1[0];
  /* dcache.vhdl:1199:34  */
  assign n24759_o = n24758_o | use_forward_rl;
  /* dcache.vhdl:1200:37  */
  assign n24760_o = r1[336];
  /* dcache.vhdl:1200:32  */
  assign n24762_o = {1'b0, n24760_o};
  /* dcache.vhdl:1201:63  */
  assign n24763_o = r1[129];
  /* dcache.vhdl:1201:44  */
  assign n24764_o = use_forward_st & n24763_o;
  /* dcache.vhdl:1203:60  */
  assign n24765_o = r1[258];
  /* dcache.vhdl:1203:42  */
  assign n24766_o = use_forward2 & n24765_o;
  /* dcache.vhdl:1203:17  */
  assign n24769_o = n24766_o ? 2'b10 : 2'b11;
  /* dcache.vhdl:1201:17  */
  assign n24771_o = n24764_o ? 2'b01 : n24769_o;
  /* dcache.vhdl:1199:17  */
  assign n24772_o = n24759_o ? n24762_o : n24771_o;
  /* dcache.vhdl:1211:68  */
  assign n24773_o = n23747_o[23:16];
  /* dcache.vhdl:1210:21  */
  assign n24775_o = n24772_o == 2'b00;
  /* dcache.vhdl:1213:64  */
  assign n24776_o = r1[86:79];
  /* dcache.vhdl:1212:21  */
  assign n24778_o = n24772_o == 2'b01;
  /* dcache.vhdl:1215:68  */
  assign n24779_o = r1[167:160];
  /* dcache.vhdl:1214:21  */
  assign n24781_o = n24772_o == 2'b10;
  /* dcache.vhdl:1217:75  */
  assign n24782_o = cache_out[23:16];
  assign n24783_o = {n24781_o, n24778_o, n24775_o};
  /* dcache.vhdl:1209:17  */
  always @*
    case (n24783_o)
      3'b100: n24784_o = n24779_o;
      3'b010: n24784_o = n24776_o;
      3'b001: n24784_o = n24773_o;
      default: n24784_o = n24782_o;
    endcase
  /* dcache.vhdl:1199:23  */
  assign n24785_o = r1[0];
  /* dcache.vhdl:1199:34  */
  assign n24786_o = n24785_o | use_forward_rl;
  /* dcache.vhdl:1200:37  */
  assign n24787_o = r1[336];
  /* dcache.vhdl:1200:32  */
  assign n24789_o = {1'b0, n24787_o};
  /* dcache.vhdl:1201:63  */
  assign n24790_o = r1[130];
  /* dcache.vhdl:1201:44  */
  assign n24791_o = use_forward_st & n24790_o;
  /* dcache.vhdl:1203:60  */
  assign n24792_o = r1[259];
  /* dcache.vhdl:1203:42  */
  assign n24793_o = use_forward2 & n24792_o;
  /* dcache.vhdl:1203:17  */
  assign n24796_o = n24793_o ? 2'b10 : 2'b11;
  /* dcache.vhdl:1201:17  */
  assign n24798_o = n24791_o ? 2'b01 : n24796_o;
  /* dcache.vhdl:1199:17  */
  assign n24799_o = n24786_o ? n24789_o : n24798_o;
  /* dcache.vhdl:1211:68  */
  assign n24800_o = n23747_o[31:24];
  /* dcache.vhdl:1210:21  */
  assign n24802_o = n24799_o == 2'b00;
  /* dcache.vhdl:1213:64  */
  assign n24803_o = r1[94:87];
  /* dcache.vhdl:1212:21  */
  assign n24805_o = n24799_o == 2'b01;
  /* dcache.vhdl:1215:68  */
  assign n24806_o = r1[175:168];
  /* dcache.vhdl:1214:21  */
  assign n24808_o = n24799_o == 2'b10;
  /* dcache.vhdl:1217:75  */
  assign n24809_o = cache_out[31:24];
  assign n24810_o = {n24808_o, n24805_o, n24802_o};
  /* dcache.vhdl:1209:17  */
  always @*
    case (n24810_o)
      3'b100: n24811_o = n24806_o;
      3'b010: n24811_o = n24803_o;
      3'b001: n24811_o = n24800_o;
      default: n24811_o = n24809_o;
    endcase
  /* dcache.vhdl:1199:23  */
  assign n24812_o = r1[0];
  /* dcache.vhdl:1199:34  */
  assign n24813_o = n24812_o | use_forward_rl;
  /* dcache.vhdl:1200:37  */
  assign n24814_o = r1[336];
  /* dcache.vhdl:1200:32  */
  assign n24816_o = {1'b0, n24814_o};
  /* dcache.vhdl:1201:63  */
  assign n24817_o = r1[131];
  /* dcache.vhdl:1201:44  */
  assign n24818_o = use_forward_st & n24817_o;
  /* dcache.vhdl:1203:60  */
  assign n24819_o = r1[260];
  /* dcache.vhdl:1203:42  */
  assign n24820_o = use_forward2 & n24819_o;
  /* dcache.vhdl:1203:17  */
  assign n24823_o = n24820_o ? 2'b10 : 2'b11;
  /* dcache.vhdl:1201:17  */
  assign n24825_o = n24818_o ? 2'b01 : n24823_o;
  /* dcache.vhdl:1199:17  */
  assign n24826_o = n24813_o ? n24816_o : n24825_o;
  /* dcache.vhdl:1211:68  */
  assign n24827_o = n23747_o[39:32];
  /* dcache.vhdl:1210:21  */
  assign n24829_o = n24826_o == 2'b00;
  /* dcache.vhdl:1213:64  */
  assign n24830_o = r1[102:95];
  /* dcache.vhdl:1212:21  */
  assign n24832_o = n24826_o == 2'b01;
  /* dcache.vhdl:1215:68  */
  assign n24833_o = r1[183:176];
  /* dcache.vhdl:1214:21  */
  assign n24835_o = n24826_o == 2'b10;
  /* dcache.vhdl:1217:75  */
  assign n24836_o = cache_out[39:32];
  assign n24837_o = {n24835_o, n24832_o, n24829_o};
  /* dcache.vhdl:1209:17  */
  always @*
    case (n24837_o)
      3'b100: n24838_o = n24833_o;
      3'b010: n24838_o = n24830_o;
      3'b001: n24838_o = n24827_o;
      default: n24838_o = n24836_o;
    endcase
  /* dcache.vhdl:1199:23  */
  assign n24839_o = r1[0];
  /* dcache.vhdl:1199:34  */
  assign n24840_o = n24839_o | use_forward_rl;
  /* dcache.vhdl:1200:37  */
  assign n24841_o = r1[336];
  /* dcache.vhdl:1200:32  */
  assign n24843_o = {1'b0, n24841_o};
  /* dcache.vhdl:1201:63  */
  assign n24844_o = r1[132];
  /* dcache.vhdl:1201:44  */
  assign n24845_o = use_forward_st & n24844_o;
  /* dcache.vhdl:1203:60  */
  assign n24846_o = r1[261];
  /* dcache.vhdl:1203:42  */
  assign n24847_o = use_forward2 & n24846_o;
  /* dcache.vhdl:1203:17  */
  assign n24850_o = n24847_o ? 2'b10 : 2'b11;
  /* dcache.vhdl:1201:17  */
  assign n24852_o = n24845_o ? 2'b01 : n24850_o;
  /* dcache.vhdl:1199:17  */
  assign n24853_o = n24840_o ? n24843_o : n24852_o;
  /* dcache.vhdl:1211:68  */
  assign n24854_o = n23747_o[47:40];
  /* dcache.vhdl:1210:21  */
  assign n24856_o = n24853_o == 2'b00;
  /* dcache.vhdl:1213:64  */
  assign n24857_o = r1[110:103];
  /* dcache.vhdl:1212:21  */
  assign n24859_o = n24853_o == 2'b01;
  /* dcache.vhdl:1215:68  */
  assign n24860_o = r1[191:184];
  /* dcache.vhdl:1214:21  */
  assign n24862_o = n24853_o == 2'b10;
  /* dcache.vhdl:1217:75  */
  assign n24863_o = cache_out[47:40];
  assign n24864_o = {n24862_o, n24859_o, n24856_o};
  /* dcache.vhdl:1209:17  */
  always @*
    case (n24864_o)
      3'b100: n24865_o = n24860_o;
      3'b010: n24865_o = n24857_o;
      3'b001: n24865_o = n24854_o;
      default: n24865_o = n24863_o;
    endcase
  /* dcache.vhdl:1199:23  */
  assign n24866_o = r1[0];
  /* dcache.vhdl:1199:34  */
  assign n24867_o = n24866_o | use_forward_rl;
  /* dcache.vhdl:1200:37  */
  assign n24868_o = r1[336];
  /* dcache.vhdl:1200:32  */
  assign n24870_o = {1'b0, n24868_o};
  /* dcache.vhdl:1201:63  */
  assign n24871_o = r1[133];
  /* dcache.vhdl:1201:44  */
  assign n24872_o = use_forward_st & n24871_o;
  /* dcache.vhdl:1203:60  */
  assign n24873_o = r1[262];
  /* dcache.vhdl:1203:42  */
  assign n24874_o = use_forward2 & n24873_o;
  /* dcache.vhdl:1203:17  */
  assign n24877_o = n24874_o ? 2'b10 : 2'b11;
  /* dcache.vhdl:1201:17  */
  assign n24879_o = n24872_o ? 2'b01 : n24877_o;
  /* dcache.vhdl:1199:17  */
  assign n24880_o = n24867_o ? n24870_o : n24879_o;
  /* dcache.vhdl:1211:68  */
  assign n24881_o = n23747_o[55:48];
  /* dcache.vhdl:1210:21  */
  assign n24883_o = n24880_o == 2'b00;
  /* dcache.vhdl:1213:64  */
  assign n24884_o = r1[118:111];
  /* dcache.vhdl:1212:21  */
  assign n24886_o = n24880_o == 2'b01;
  /* dcache.vhdl:1215:68  */
  assign n24887_o = r1[199:192];
  /* dcache.vhdl:1214:21  */
  assign n24889_o = n24880_o == 2'b10;
  /* dcache.vhdl:1217:75  */
  assign n24890_o = cache_out[55:48];
  assign n24891_o = {n24889_o, n24886_o, n24883_o};
  /* dcache.vhdl:1209:17  */
  always @*
    case (n24891_o)
      3'b100: n24892_o = n24887_o;
      3'b010: n24892_o = n24884_o;
      3'b001: n24892_o = n24881_o;
      default: n24892_o = n24890_o;
    endcase
  /* dcache.vhdl:1199:23  */
  assign n24893_o = r1[0];
  /* dcache.vhdl:1199:34  */
  assign n24894_o = n24893_o | use_forward_rl;
  /* dcache.vhdl:1200:37  */
  assign n24895_o = r1[336];
  /* dcache.vhdl:1200:32  */
  assign n24897_o = {1'b0, n24895_o};
  /* dcache.vhdl:1201:63  */
  assign n24898_o = r1[134];
  /* dcache.vhdl:1201:44  */
  assign n24899_o = use_forward_st & n24898_o;
  /* dcache.vhdl:1203:60  */
  assign n24900_o = r1[263];
  /* dcache.vhdl:1203:42  */
  assign n24901_o = use_forward2 & n24900_o;
  /* dcache.vhdl:1203:17  */
  assign n24904_o = n24901_o ? 2'b10 : 2'b11;
  /* dcache.vhdl:1201:17  */
  assign n24906_o = n24899_o ? 2'b01 : n24904_o;
  /* dcache.vhdl:1199:17  */
  assign n24907_o = n24894_o ? n24897_o : n24906_o;
  /* dcache.vhdl:1211:68  */
  assign n24908_o = n23747_o[63:56];
  /* dcache.vhdl:1210:21  */
  assign n24910_o = n24907_o == 2'b00;
  /* dcache.vhdl:1213:64  */
  assign n24911_o = r1[126:119];
  /* dcache.vhdl:1212:21  */
  assign n24913_o = n24907_o == 2'b01;
  /* dcache.vhdl:1215:68  */
  assign n24914_o = r1[207:200];
  /* dcache.vhdl:1214:21  */
  assign n24916_o = n24907_o == 2'b10;
  /* dcache.vhdl:1217:75  */
  assign n24917_o = cache_out[63:56];
  assign n24918_o = {n24916_o, n24913_o, n24910_o};
  /* dcache.vhdl:1209:17  */
  always @*
    case (n24918_o)
      3'b100: n24919_o = n24914_o;
      3'b010: n24919_o = n24911_o;
      3'b001: n24919_o = n24908_o;
      default: n24919_o = n24917_o;
    endcase
  assign n24920_o = {n24919_o, n24892_o, n24865_o, n24838_o, n24811_o, n24784_o, n24757_o, n24730_o};
  /* dcache.vhdl:1223:34  */
  assign n24921_o = r1[491:444];
  /* dcache.vhdl:1224:34  */
  assign n24922_o = r1[496:492];
  /* dcache.vhdl:1226:36  */
  assign n24923_o = r1[337];
  /* dcache.vhdl:1227:19  */
  assign n24924_o = r1[335:334];
  /* dcache.vhdl:1227:25  */
  assign n24926_o = n24924_o == 2'b01;
  /* dcache.vhdl:1227:59  */
  assign n24927_o = n23747_o[64];
  /* dcache.vhdl:1227:43  */
  assign n24928_o = n24926_o & n24927_o;
  /* dcache.vhdl:1227:13  */
  assign n24930_o = n24928_o ? 1'b1 : n24923_o;
  /* dcache.vhdl:1234:23  */
  assign n24932_o = req_op == 3'b011;
  /* dcache.vhdl:1234:13  */
  assign n24935_o = n24932_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:1239:23  */
  assign n24937_o = req_op == 3'b011;
  /* dcache.vhdl:1239:47  */
  assign n24939_o = req_op == 3'b110;
  /* dcache.vhdl:1239:37  */
  assign n24940_o = n24937_o | n24939_o;
  /* dcache.vhdl:1239:13  */
  assign n24943_o = n24940_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:1245:23  */
  assign n24945_o = req_op == 3'b001;
  /* dcache.vhdl:1248:39  */
  assign n24946_o = r0[149];
  /* dcache.vhdl:1248:32  */
  assign n24947_o = ~n24946_o;
  /* dcache.vhdl:1249:36  */
  assign n24948_o = r0[149];
  assign n24952_o = {1'b0, 1'b0};
  assign n24953_o = {access_ok, n24948_o};
  /* dcache.vhdl:1245:13  */
  assign n24954_o = n24945_o ? n24947_o : 1'b0;
  /* dcache.vhdl:1245:13  */
  assign n24955_o = n24945_o ? n24953_o : n24952_o;
  /* dcache.vhdl:1257:23  */
  assign n24957_o = req_op == 3'b010;
  /* dcache.vhdl:1257:13  */
  assign n24960_o = n24957_o ? 1'b1 : 1'b0;
  assign n24961_o = {n24920_o, n24922_o, n24930_o, ram_wr_select, n24921_o, ram_wr_data, tlb_req_index, tlb_hit_way, tlb_hit, n24943_o, req_index, n24935_o};
  assign n24962_o = {n24960_o, n24955_o};
  /* dcache.vhdl:1316:49  */
  assign n25002_o = r0[146];
  /* dcache.vhdl:1316:61  */
  assign n25003_o = r0[148];
  /* dcache.vhdl:1316:55  */
  assign n25004_o = n25002_o | n25003_o;
  /* dcache.vhdl:1316:41  */
  assign n25005_o = r0_valid & n25004_o;
  /* dcache.vhdl:1317:27  */
  assign n25007_o = req_op == 3'b011;
  /* dcache.vhdl:1317:51  */
  assign n25009_o = req_op == 3'b010;
  /* dcache.vhdl:1317:41  */
  assign n25010_o = n25007_o | n25009_o;
  /* dcache.vhdl:1318:27  */
  assign n25011_o = r0[149];
  /* dcache.vhdl:1318:35  */
  assign n25012_o = ~n25011_o;
  /* dcache.vhdl:1317:17  */
  assign n25015_o = n25017_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:1318:21  */
  assign n25016_o = n25012_o ? n25005_o : 1'b1;
  /* dcache.vhdl:1317:17  */
  assign n25017_o = n25010_o & n25012_o;
  /* dcache.vhdl:1317:17  */
  assign n25018_o = n25010_o ? n25016_o : n25005_o;
  /* dcache.vhdl:1327:73  */
  assign n25024_o = snoop_tag_set == snoop_wrtag;
  /* dcache.vhdl:1327:42  */
  assign n25025_o = snoop_valid & n25024_o;
  /* dcache.vhdl:1328:38  */
  assign n25027_o = 2'b11 - snoop_index;
  /* dcache.vhdl:1327:21  */
  assign n25031_o = n25025_o ? n25919_o : cache_valids;
  /* dcache.vhdl:1332:23  */
  assign n25032_o = r1[338];
  /* dcache.vhdl:1336:43  */
  assign n25033_o = r1[498:497];
  /* dcache.vhdl:1337:72  */
  assign n25037_o = r1[491:444];
  assign n25042_o = r1[338];
  /* dcache.vhdl:1332:17  */
  assign n25043_o = n25032_o ? 1'b0 : n25042_o;
  /* dcache.vhdl:1346:23  */
  assign n25044_o = r1[0];
  /* dcache.vhdl:1347:31  */
  assign n25045_o = r1[136:2];
  /* dcache.vhdl:1351:39  */
  assign n25046_o = r0[149];
  /* dcache.vhdl:1352:36  */
  assign n25047_o = r0[145:0];
  /* dcache.vhdl:1352:40  */
  assign n25048_o = n25047_o[3];
  /* dcache.vhdl:1355:27  */
  assign n25049_o = r0[145:0];
  /* dcache.vhdl:1355:31  */
  assign n25050_o = n25049_o[3];
  /* dcache.vhdl:1357:30  */
  assign n25052_o = r0[150];
  /* dcache.vhdl:1358:40  */
  assign n25053_o = r0[145:0];
  /* dcache.vhdl:1358:44  */
  assign n25054_o = n25053_o[137:74];
  /* dcache.vhdl:1360:42  */
  assign n25055_o = n23725_o[137:74];
  /* dcache.vhdl:1357:21  */
  assign n25056_o = n25052_o ? n25054_o : n25055_o;
  /* dcache.vhdl:1355:21  */
  assign n25057_o = n25050_o ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n25056_o;
  /* dcache.vhdl:1363:27  */
  assign n25058_o = r0[145:0];
  /* dcache.vhdl:1363:31  */
  assign n25059_o = n25058_o[3];
  /* dcache.vhdl:1363:49  */
  assign n25060_o = r0[145:0];
  /* dcache.vhdl:1363:53  */
  assign n25061_o = n25060_o[2];
  /* dcache.vhdl:1363:71  */
  assign n25062_o = r0[145:0];
  /* dcache.vhdl:1363:75  */
  assign n25063_o = n25062_o[4];
  /* dcache.vhdl:1363:78  */
  assign n25064_o = ~n25063_o;
  /* dcache.vhdl:1363:64  */
  assign n25065_o = n25061_o & n25064_o;
  /* dcache.vhdl:1363:98  */
  assign n25066_o = perm_attr[2];
  /* dcache.vhdl:1363:106  */
  assign n25067_o = ~n25066_o;
  /* dcache.vhdl:1363:84  */
  assign n25068_o = n25065_o & n25067_o;
  /* dcache.vhdl:1363:42  */
  assign n25069_o = n25059_o | n25068_o;
  /* dcache.vhdl:1366:44  */
  assign n25071_o = r0[145:0];
  /* dcache.vhdl:1366:48  */
  assign n25072_o = n25071_o[145:138];
  /* dcache.vhdl:1363:21  */
  assign n25073_o = n25069_o ? 8'b11111111 : n25072_o;
  /* dcache.vhdl:1373:31  */
  assign n25075_o = req_op == 3'b100;
  /* dcache.vhdl:1373:56  */
  assign n25077_o = req_op == 3'b101;
  /* dcache.vhdl:1373:46  */
  assign n25078_o = n25075_o | n25077_o;
  /* dcache.vhdl:1374:32  */
  assign n25080_o = req_op == 3'b111;
  /* dcache.vhdl:1373:69  */
  assign n25081_o = n25078_o | n25080_o;
  /* dcache.vhdl:1374:58  */
  assign n25083_o = req_op == 3'b110;
  /* dcache.vhdl:1374:48  */
  assign n25084_o = n25081_o | n25083_o;
  assign n25085_o = {n25046_o, req_same_tag, n25073_o, n25057_o, ra, n25048_o, req_go, req_op};
  assign n25087_o = r1[0];
  /* dcache.vhdl:1373:21  */
  assign n25088_o = n25084_o ? 1'b1 : n25087_o;
  assign n25091_o = r1[0];
  /* dcache.vhdl:1346:17  */
  assign n25092_o = n25044_o ? n25091_o : n25088_o;
  assign n25095_o = {n25046_o, req_same_tag, n25073_o, n25057_o, ra, n25048_o, req_go, req_op};
  /* dcache.vhdl:1346:17  */
  assign n25096_o = n25044_o ? n25045_o : n25095_o;
  /* dcache.vhdl:1381:25  */
  assign n25097_o = r1[335:334];
  /* dcache.vhdl:1383:49  */
  assign n25099_o = n25096_o[60:5];
  /* wishbone_types.vhdl:69:20  */
  assign n25104_o = n25099_o[31:3];
  /* dcache.vhdl:1384:38  */
  assign n25105_o = n25096_o[132:125];
  /* dcache.vhdl:1385:38  */
  assign n25106_o = n25096_o[124:61];
  /* dcache.vhdl:1386:36  */
  assign n25107_o = n25096_o[4];
  /* dcache.vhdl:1389:53  */
  assign n25109_o = n25096_o[60:5];
  /* dcache.vhdl:437:40  */
  assign n25114_o = n25109_o[7:6];
  /* dcache.vhdl:1390:49  */
  assign n25117_o = n25096_o[60:5];
  /* dcache.vhdl:443:40  */
  assign n25122_o = n25117_o[7:3];
  /* dcache.vhdl:1391:66  */
  assign n25126_o = n25096_o[60:5];
  /* dcache.vhdl:443:40  */
  assign n25131_o = n25126_o[7:3];
  /* dcache.vhdl:451:21  */
  assign n25140_o = n25131_o[2:0];
  /* dcache.vhdl:1391:78  */
  assign n25142_o = n25140_o - 3'b001;
  /* dcache.vhdl:1392:50  */
  assign n25144_o = n25096_o[60:5];
  /* dcache.vhdl:497:20  */
  assign n25149_o = n25144_o[55:8];
  /* dcache.vhdl:1404:30  */
  assign n25162_o = n25096_o[2:0];
  /* dcache.vhdl:1405:21  */
  assign n25164_o = n25162_o == 3'b011;
  /* dcache.vhdl:1408:21  */
  assign n25172_o = n25162_o == 3'b100;
  /* dcache.vhdl:1425:21  */
  assign n25178_o = n25162_o == 3'b101;
  /* dcache.vhdl:1432:32  */
  assign n25179_o = n25096_o[4];
  /* dcache.vhdl:1432:37  */
  assign n25180_o = ~n25179_o;
  /* dcache.vhdl:1437:36  */
  assign n25185_o = n25096_o[134];
  /* dcache.vhdl:1437:44  */
  assign n25186_o = ~n25185_o;
  /* dcache.vhdl:1432:25  */
  assign n25189_o = n25209_o ? 1'b1 : n25015_o;
  /* dcache.vhdl:1437:29  */
  assign n25190_o = n25186_o ? n25018_o : 1'b1;
  /* dcache.vhdl:1442:36  */
  assign n25191_o = n25096_o[2:0];
  /* dcache.vhdl:1442:39  */
  assign n25193_o = n25191_o == 3'b110;
  /* dcache.vhdl:1432:25  */
  assign n25195_o = n25204_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:1449:36  */
  assign n25197_o = n25096_o[2:0];
  /* dcache.vhdl:1449:39  */
  assign n25199_o = n25197_o == 3'b111;
  /* dcache.vhdl:1449:29  */
  assign n25201_o = n25199_o ? 1'b1 : n25043_o;
  /* dcache.vhdl:1432:25  */
  assign n25202_o = n25180_o ? 1'b0 : n25092_o;
  /* dcache.vhdl:1432:25  */
  assign n25203_o = n25180_o ? 2'b10 : 2'b01;
  /* dcache.vhdl:1432:25  */
  assign n25204_o = n25180_o & n25193_o;
  /* dcache.vhdl:1432:25  */
  assign n25205_o = n25180_o ? n25043_o : n25201_o;
  /* dcache.vhdl:1432:25  */
  assign n25206_o = n25180_o ? 1'b1 : 1'b0;
  assign n25207_o = r1[512:510];
  /* dcache.vhdl:1432:25  */
  assign n25208_o = n25180_o ? 3'b001 : n25207_o;
  /* dcache.vhdl:1432:25  */
  assign n25209_o = n25180_o & n25186_o;
  /* dcache.vhdl:1432:25  */
  assign n25210_o = n25180_o ? n25190_o : n25018_o;
  /* dcache.vhdl:1456:32  */
  assign n25214_o = n25096_o[2:0];
  /* dcache.vhdl:1456:35  */
  assign n25216_o = n25214_o == 3'b111;
  /* dcache.vhdl:1456:25  */
  assign n25218_o = n25216_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:1431:21  */
  assign n25220_o = n25162_o == 3'b110;
  /* dcache.vhdl:1431:39  */
  assign n25222_o = n25162_o == 3'b111;
  /* dcache.vhdl:1431:39  */
  assign n25223_o = n25220_o | n25222_o;
  /* dcache.vhdl:1462:21  */
  assign n25225_o = n25162_o == 3'b000;
  /* dcache.vhdl:1463:21  */
  assign n25227_o = n25162_o == 3'b001;
  /* dcache.vhdl:1464:21  */
  assign n25229_o = n25162_o == 3'b010;
  assign n25230_o = {n25229_o, n25227_o, n25225_o, n25223_o, n25178_o, n25172_o, n25164_o};
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25232_o = n25092_o;
      7'b0100000: n25232_o = n25092_o;
      7'b0010000: n25232_o = n25092_o;
      7'b0001000: n25232_o = n25202_o;
      7'b0000100: n25232_o = n25092_o;
      7'b0000010: n25232_o = n25092_o;
      7'b0000001: n25232_o = n25092_o;
      default: n25232_o = 1'bX;
    endcase
  assign n25233_o = r1[335:334];
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25235_o = n25233_o;
      7'b0100000: n25235_o = n25233_o;
      7'b0010000: n25235_o = n25233_o;
      7'b0001000: n25235_o = n25203_o;
      7'b0000100: n25235_o = 2'b11;
      7'b0000010: n25235_o = 2'b01;
      7'b0000001: n25235_o = n25233_o;
      default: n25235_o = 2'bX;
    endcase
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25237_o = 1'b0;
      7'b0100000: n25237_o = 1'b0;
      7'b0010000: n25237_o = 1'b0;
      7'b0001000: n25237_o = n25195_o;
      7'b0000100: n25237_o = 1'b0;
      7'b0000010: n25237_o = 1'b0;
      7'b0000001: n25237_o = 1'b0;
      default: n25237_o = 1'bX;
    endcase
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25239_o = n25043_o;
      7'b0100000: n25239_o = n25043_o;
      7'b0010000: n25239_o = n25043_o;
      7'b0001000: n25239_o = n25205_o;
      7'b0000100: n25239_o = n25043_o;
      7'b0000010: n25239_o = 1'b1;
      7'b0000001: n25239_o = n25043_o;
      default: n25239_o = 1'bX;
    endcase
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25241_o = 1'b0;
      7'b0100000: n25241_o = 1'b0;
      7'b0010000: n25241_o = 1'b0;
      7'b0001000: n25241_o = n25206_o;
      7'b0000100: n25241_o = 1'b0;
      7'b0000010: n25241_o = 1'b0;
      7'b0000001: n25241_o = 1'b0;
      default: n25241_o = 1'bX;
    endcase
  assign n25242_o = r1[441];
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25244_o = n25242_o;
      7'b0100000: n25244_o = n25242_o;
      7'b0010000: n25244_o = n25242_o;
      7'b0001000: n25244_o = 1'b1;
      7'b0000100: n25244_o = 1'b1;
      7'b0000010: n25244_o = 1'b1;
      7'b0000001: n25244_o = n25242_o;
      default: n25244_o = 1'bX;
    endcase
  assign n25245_o = r1[442];
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25247_o = n25245_o;
      7'b0100000: n25247_o = n25245_o;
      7'b0010000: n25247_o = n25245_o;
      7'b0001000: n25247_o = 1'b1;
      7'b0000100: n25247_o = 1'b1;
      7'b0000010: n25247_o = 1'b1;
      7'b0000001: n25247_o = n25245_o;
      default: n25247_o = 1'bX;
    endcase
  assign n25248_o = r1[443];
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25250_o = n25248_o;
      7'b0100000: n25250_o = n25248_o;
      7'b0010000: n25250_o = n25248_o;
      7'b0001000: n25250_o = 1'b1;
      7'b0000100: n25250_o = 1'b0;
      7'b0000010: n25250_o = 1'b0;
      7'b0000001: n25250_o = n25248_o;
      default: n25250_o = 1'bX;
    endcase
  assign n25251_o = r1[512:510];
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25253_o = n25251_o;
      7'b0100000: n25253_o = n25251_o;
      7'b0010000: n25253_o = n25251_o;
      7'b0001000: n25253_o = n25208_o;
      7'b0000100: n25253_o = n25251_o;
      7'b0000010: n25253_o = n25251_o;
      7'b0000001: n25253_o = n25251_o;
      default: n25253_o = 3'bX;
    endcase
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25255_o = n25015_o;
      7'b0100000: n25255_o = n25015_o;
      7'b0010000: n25255_o = n25015_o;
      7'b0001000: n25255_o = n25189_o;
      7'b0000100: n25255_o = n25015_o;
      7'b0000010: n25255_o = n25015_o;
      7'b0000001: n25255_o = n25015_o;
      default: n25255_o = 1'bX;
    endcase
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25257_o = n25018_o;
      7'b0100000: n25257_o = n25018_o;
      7'b0010000: n25257_o = n25018_o;
      7'b0001000: n25257_o = n25210_o;
      7'b0000100: n25257_o = n25018_o;
      7'b0000010: n25257_o = n25018_o;
      7'b0000001: n25257_o = n25018_o;
      default: n25257_o = 1'bX;
    endcase
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25259_o = 1'b0;
      7'b0100000: n25259_o = 1'b0;
      7'b0010000: n25259_o = 1'b0;
      7'b0001000: n25259_o = 1'b0;
      7'b0000100: n25259_o = 1'b0;
      7'b0000010: n25259_o = 1'b1;
      7'b0000001: n25259_o = 1'b0;
      default: n25259_o = 1'bX;
    endcase
  /* dcache.vhdl:1404:21  */
  always @*
    case (n25230_o)
      7'b1000000: n25261_o = 1'b0;
      7'b0100000: n25261_o = 1'b0;
      7'b0010000: n25261_o = 1'b0;
      7'b0001000: n25261_o = n25218_o;
      7'b0000100: n25261_o = 1'b0;
      7'b0000010: n25261_o = 1'b0;
      7'b0000001: n25261_o = 1'b0;
      default: n25261_o = 1'bX;
    endcase
  /* dcache.vhdl:1382:17  */
  assign n25263_o = n25097_o == 2'b00;
  /* dcache.vhdl:1469:36  */
  assign n25264_o = n23747_o[65];
  /* dcache.vhdl:1469:42  */
  assign n25265_o = ~n25264_o;
  /* dcache.vhdl:1469:55  */
  assign n25266_o = r1[443:340];
  /* dcache.vhdl:1469:58  */
  assign n25267_o = n25266_o[102];
  /* dcache.vhdl:1469:48  */
  assign n25268_o = n25265_o & n25267_o;
  /* dcache.vhdl:1471:51  */
  assign n25270_o = r1[443:340];
  /* dcache.vhdl:1471:54  */
  assign n25271_o = n25270_o[28:0];
  /* dcache.vhdl:1471:62  */
  assign n25272_o = r1[501:499];
  /* dcache.vhdl:457:29  */
  assign n25277_o = n25271_o[2:0];
  /* dcache.vhdl:457:74  */
  assign n25278_o = n25277_o == n25272_o;
  assign n25280_o = r1[442];
  /* dcache.vhdl:1469:21  */
  assign n25281_o = n25301_o ? 1'b0 : n25280_o;
  /* dcache.vhdl:1476:58  */
  assign n25283_o = r1[443:340];
  /* dcache.vhdl:1476:61  */
  assign n25284_o = n25283_o[28:0];
  /* dcache.vhdl:472:24  */
  assign n25291_o = n25284_o[2:0];
  /* dcache.vhdl:473:56  */
  assign n25294_o = n25291_o + 3'b001;
  assign n25296_o = r1[368:343];
  assign n25297_o = {n25296_o, n25294_o};
  assign n25298_o = r1[368:340];
  /* dcache.vhdl:1469:21  */
  assign n25299_o = n25268_o ? n25297_o : n25298_o;
  /* dcache.vhdl:1469:21  */
  assign n25301_o = n25268_o & n25278_o;
  /* dcache.vhdl:1480:36  */
  assign n25302_o = n23747_o[64];
  /* dcache.vhdl:1481:42  */
  assign n25303_o = r1[496:492];
  /* dcache.vhdl:1481:52  */
  assign n25304_o = {27'b0, n25303_o};  //  uext
  assign n25305_o = n25304_o[2:0];
  /* dcache.vhdl:1481:52  */
  assign n25308_o = 3'b111 - n25305_o;
  assign n25310_o = r1[509:502];
  /* dcache.vhdl:1488:31  */
  assign n25313_o = r1[0];
  /* dcache.vhdl:1488:49  */
  assign n25314_o = r1[136:2];
  /* dcache.vhdl:1488:53  */
  assign n25315_o = n25314_o[133];
  /* dcache.vhdl:1488:42  */
  assign n25316_o = n25313_o & n25315_o;
  /* dcache.vhdl:1489:34  */
  assign n25317_o = r1[336];
  /* dcache.vhdl:1489:53  */
  assign n25318_o = n25096_o[4];
  /* dcache.vhdl:1489:45  */
  assign n25319_o = n25317_o & n25318_o;
  /* dcache.vhdl:1489:71  */
  assign n25320_o = r1[136:2];
  /* dcache.vhdl:1489:75  */
  assign n25321_o = n25320_o[2:0];
  /* dcache.vhdl:1489:78  */
  assign n25323_o = n25321_o == 3'b100;
  /* dcache.vhdl:1489:65  */
  assign n25324_o = n25319_o | n25323_o;
  /* dcache.vhdl:1488:68  */
  assign n25325_o = n25316_o & n25324_o;
  /* dcache.vhdl:1490:32  */
  assign n25326_o = r1[496:492];
  /* dcache.vhdl:1490:42  */
  assign n25327_o = {27'b0, n25326_o};  //  uext
  /* dcache.vhdl:1490:55  */
  assign n25329_o = r1[136:2];
  /* dcache.vhdl:1490:59  */
  assign n25330_o = n25329_o[60:5];
  /* dcache.vhdl:443:40  */
  assign n25335_o = n25330_o[7:3];
  /* dcache.vhdl:1490:42  */
  assign n25337_o = {27'b0, n25335_o};  //  uext
  /* dcache.vhdl:1490:42  */
  assign n25338_o = n25327_o == n25337_o;
  /* dcache.vhdl:1489:94  */
  assign n25339_o = n25325_o & n25338_o;
  /* dcache.vhdl:1493:35  */
  assign n25342_o = r1[1];
  /* dcache.vhdl:1493:43  */
  assign n25343_o = ~n25342_o;
  /* dcache.vhdl:1480:21  */
  assign n25346_o = n25414_o ? 1'b1 : n25015_o;
  /* dcache.vhdl:1493:29  */
  assign n25347_o = n25343_o ? n25018_o : 1'b1;
  /* dcache.vhdl:1480:21  */
  assign n25348_o = n25404_o ? 1'b0 : n25092_o;
  /* dcache.vhdl:1480:21  */
  assign n25349_o = n25407_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:1488:25  */
  assign n25350_o = n25339_o & n25343_o;
  /* dcache.vhdl:1480:21  */
  assign n25351_o = n25415_o ? n25347_o : n25018_o;
  /* dcache.vhdl:1501:43  */
  assign n25353_o = r1[496:492];
  /* dcache.vhdl:1501:57  */
  assign n25354_o = r1[501:499];
  /* dcache.vhdl:451:21  */
  assign n25367_o = n25353_o[2:0];
  /* dcache.vhdl:463:37  */
  assign n25368_o = n25367_o == n25354_o;
  /* dcache.vhdl:1506:45  */
  assign n25370_o = r1[498:497];
  /* dcache.vhdl:1506:45  */
  assign n25372_o = 2'b11 - n25370_o;
  /* dcache.vhdl:1508:56  */
  assign n25376_o = r1[336];
  /* dcache.vhdl:1508:49  */
  assign n25377_o = ~n25376_o;
  /* dcache.vhdl:1480:21  */
  assign n25379_o = n25403_o ? n25971_o : n25031_o;
  assign n25380_o = r1[335:334];
  /* dcache.vhdl:1480:21  */
  assign n25381_o = n25406_o ? 2'b00 : n25380_o;
  assign n25382_o = r1[441];
  /* dcache.vhdl:1480:21  */
  assign n25383_o = n25409_o ? 1'b0 : n25382_o;
  /* dcache.vhdl:1480:21  */
  assign n25384_o = n25416_o ? n25377_o : 1'b0;
  /* dcache.vhdl:1513:53  */
  assign n25386_o = r1[496:492];
  /* dcache.vhdl:489:24  */
  assign n25396_o = n25386_o[2:0];
  /* dcache.vhdl:490:78  */
  assign n25399_o = n25396_o + 3'b001;
  assign n25400_o = r1[496:495];
  assign n25401_o = {n25400_o, n25399_o};
  /* dcache.vhdl:1480:21  */
  assign n25403_o = n25302_o & n25368_o;
  /* dcache.vhdl:1480:21  */
  assign n25404_o = n25302_o & n25339_o;
  /* dcache.vhdl:1480:21  */
  assign n25406_o = n25302_o & n25368_o;
  /* dcache.vhdl:1480:21  */
  assign n25407_o = n25302_o & n25339_o;
  /* dcache.vhdl:1480:21  */
  assign n25409_o = n25302_o & n25368_o;
  assign n25410_o = r1[496:492];
  /* dcache.vhdl:1480:21  */
  assign n25411_o = n25302_o ? n25401_o : n25410_o;
  assign n25412_o = r1[509:502];
  /* dcache.vhdl:1480:21  */
  assign n25413_o = n25302_o ? n25954_o : n25412_o;
  /* dcache.vhdl:1480:21  */
  assign n25414_o = n25302_o & n25350_o;
  /* dcache.vhdl:1480:21  */
  assign n25415_o = n25302_o & n25339_o;
  /* dcache.vhdl:1480:21  */
  assign n25416_o = n25302_o & n25368_o;
  /* dcache.vhdl:1467:17  */
  assign n25418_o = n25097_o == 2'b01;
  /* dcache.vhdl:1517:37  */
  assign n25419_o = r1[443:340];
  /* dcache.vhdl:1517:40  */
  assign n25420_o = n25419_o[102];
  /* dcache.vhdl:1517:44  */
  assign n25421_o = ~n25420_o;
  /* dcache.vhdl:1518:32  */
  assign n25422_o = r1[512:510];
  /* dcache.vhdl:1519:27  */
  assign n25423_o = r1[513];
  /* dcache.vhdl:1519:42  */
  assign n25424_o = r1[514];
  /* dcache.vhdl:1519:36  */
  assign n25425_o = n25423_o != n25424_o;
  /* dcache.vhdl:1520:31  */
  assign n25426_o = r1[513];
  /* dcache.vhdl:1521:42  */
  assign n25428_o = n25422_o + 3'b001;
  /* dcache.vhdl:1523:42  */
  assign n25430_o = n25422_o - 3'b001;
  /* dcache.vhdl:1520:25  */
  assign n25431_o = n25426_o ? n25428_o : n25430_o;
  /* dcache.vhdl:1519:21  */
  assign n25432_o = n25425_o ? n25431_o : n25422_o;
  /* dcache.vhdl:1528:36  */
  assign n25433_o = n23747_o[65];
  /* dcache.vhdl:1528:42  */
  assign n25434_o = ~n25433_o;
  /* dcache.vhdl:1531:32  */
  assign n25435_o = n25096_o[3];
  /* dcache.vhdl:1533:46  */
  assign n25436_o = n25096_o[12:8];
  /* dcache.vhdl:1534:46  */
  assign n25437_o = n25096_o[124:61];
  /* dcache.vhdl:1535:46  */
  assign n25438_o = n25096_o[132:125];
  assign n25439_o = {n25438_o, n25437_o};
  assign n25440_o = r1[344:340];
  /* dcache.vhdl:1531:25  */
  assign n25441_o = n25435_o ? n25436_o : n25440_o;
  assign n25442_o = r1[440:369];
  /* dcache.vhdl:1528:21  */
  assign n25443_o = n25496_o ? n25439_o : n25442_o;
  /* dcache.vhdl:1537:33  */
  assign n25445_o = $unsigned(n25432_o) < $unsigned(3'b111);
  /* dcache.vhdl:1537:45  */
  assign n25446_o = n25096_o[133];
  /* dcache.vhdl:1537:37  */
  assign n25447_o = n25445_o & n25446_o;
  /* dcache.vhdl:1537:68  */
  assign n25448_o = n25096_o[4];
  /* dcache.vhdl:1537:73  */
  assign n25449_o = ~n25448_o;
  /* dcache.vhdl:1537:60  */
  assign n25450_o = n25447_o & n25449_o;
  /* dcache.vhdl:1538:34  */
  assign n25451_o = n25096_o[2:0];
  /* dcache.vhdl:1538:37  */
  assign n25453_o = n25451_o == 3'b111;
  /* dcache.vhdl:1538:60  */
  assign n25454_o = n25096_o[2:0];
  /* dcache.vhdl:1538:63  */
  assign n25456_o = n25454_o == 3'b110;
  /* dcache.vhdl:1538:53  */
  assign n25457_o = n25453_o | n25456_o;
  /* dcache.vhdl:1537:79  */
  assign n25458_o = n25450_o & n25457_o;
  /* dcache.vhdl:1542:57  */
  assign n25461_o = n25096_o[60:5];
  /* dcache.vhdl:443:40  */
  assign n25466_o = n25461_o[7:3];
  /* dcache.vhdl:1543:36  */
  assign n25468_o = n25096_o[2:0];
  /* dcache.vhdl:1543:39  */
  assign n25470_o = n25468_o == 3'b110;
  /* dcache.vhdl:1528:21  */
  assign n25472_o = n25491_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:1528:21  */
  assign n25478_o = n25490_o ? 1'b0 : n25092_o;
  /* dcache.vhdl:1537:25  */
  assign n25479_o = n25458_o & n25470_o;
  /* dcache.vhdl:1537:25  */
  assign n25480_o = n25458_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:1537:25  */
  assign n25481_o = n25458_o ? 1'b1 : 1'b0;
  assign n25482_o = r1[496:492];
  /* dcache.vhdl:1528:21  */
  assign n25483_o = n25500_o ? n25466_o : n25482_o;
  /* dcache.vhdl:1528:21  */
  assign n25484_o = n25501_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:1528:21  */
  assign n25485_o = n25502_o ? 1'b1 : n25015_o;
  /* dcache.vhdl:1537:25  */
  assign n25488_o = n25458_o ? 1'b0 : 1'b1;
  assign n25489_o = {n25441_o, n25480_o};
  /* dcache.vhdl:1528:21  */
  assign n25490_o = n25434_o & n25458_o;
  /* dcache.vhdl:1528:21  */
  assign n25491_o = n25434_o & n25479_o;
  assign n25492_o = r1[344:340];
  assign n25493_o = {n25492_o, 1'b0};
  /* dcache.vhdl:1528:21  */
  assign n25494_o = n25434_o ? n25489_o : n25493_o;
  /* dcache.vhdl:1528:21  */
  assign n25496_o = n25434_o & n25435_o;
  assign n25497_o = r1[442];
  /* dcache.vhdl:1528:21  */
  assign n25498_o = n25434_o ? n25481_o : n25497_o;
  /* dcache.vhdl:1528:21  */
  assign n25500_o = n25434_o & n25458_o;
  /* dcache.vhdl:1528:21  */
  assign n25501_o = n25434_o & n25458_o;
  /* dcache.vhdl:1528:21  */
  assign n25502_o = n25434_o & n25458_o;
  /* dcache.vhdl:1528:21  */
  assign n25503_o = n25434_o ? n25488_o : n25421_o;
  /* dcache.vhdl:1559:36  */
  assign n25504_o = n23747_o[64];
  /* dcache.vhdl:1560:47  */
  assign n25506_o = n25432_o == 3'b001;
  /* dcache.vhdl:1560:38  */
  assign n25507_o = n25503_o & n25506_o;
  assign n25511_o = {1'b0, 1'b0};
  assign n25512_o = r1[335:334];
  /* dcache.vhdl:1559:21  */
  assign n25513_o = n25519_o ? 2'b00 : n25512_o;
  assign n25514_o = r1[441];
  assign n25515_o = {n25498_o, n25514_o};
  /* dcache.vhdl:1560:25  */
  assign n25516_o = n25507_o ? n25511_o : n25515_o;
  /* dcache.vhdl:1559:21  */
  assign n25519_o = n25504_o & n25507_o;
  assign n25520_o = r1[441];
  assign n25521_o = {n25498_o, n25520_o};
  /* dcache.vhdl:1559:21  */
  assign n25522_o = n25504_o ? n25516_o : n25521_o;
  /* dcache.vhdl:1559:21  */
  assign n25523_o = n25504_o ? 1'b1 : 1'b0;
  /* dcache.vhdl:1516:17  */
  assign n25525_o = n25097_o == 2'b10;
  /* dcache.vhdl:1570:36  */
  assign n25526_o = n23747_o[65];
  /* dcache.vhdl:1570:42  */
  assign n25527_o = ~n25526_o;
  assign n25529_o = r1[442];
  /* dcache.vhdl:1570:21  */
  assign n25530_o = n25527_o ? 1'b0 : n25529_o;
  /* dcache.vhdl:1575:36  */
  assign n25531_o = n23747_o[64];
  /* dcache.vhdl:1579:31  */
  assign n25535_o = r1[1];
  /* dcache.vhdl:1579:39  */
  assign n25536_o = ~n25535_o;
  /* dcache.vhdl:1575:21  */
  assign n25539_o = n25551_o ? 1'b1 : n25015_o;
  /* dcache.vhdl:1579:25  */
  assign n25540_o = n25536_o ? n25018_o : 1'b1;
  assign n25543_o = {1'b0, 1'b0};
  /* dcache.vhdl:1575:21  */
  assign n25544_o = n25531_o ? 1'b0 : n25092_o;
  assign n25545_o = r1[335:334];
  /* dcache.vhdl:1575:21  */
  assign n25546_o = n25531_o ? 2'b00 : n25545_o;
  /* dcache.vhdl:1575:21  */
  assign n25547_o = n25531_o ? 1'b1 : 1'b0;
  assign n25548_o = r1[441];
  assign n25549_o = {n25530_o, n25548_o};
  /* dcache.vhdl:1575:21  */
  assign n25550_o = n25531_o ? n25543_o : n25549_o;
  /* dcache.vhdl:1575:21  */
  assign n25551_o = n25531_o & n25536_o;
  /* dcache.vhdl:1575:21  */
  assign n25552_o = n25531_o ? n25540_o : n25018_o;
  /* dcache.vhdl:1568:17  */
  assign n25554_o = n25097_o == 2'b11;
  assign n25555_o = {n25554_o, n25525_o, n25418_o, n25263_o};
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25557_o = n25031_o;
      4'b0100: n25557_o = n25031_o;
      4'b0010: n25557_o = n25379_o;
      4'b0001: n25557_o = n25031_o;
      default: n25557_o = 4'bX;
    endcase
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25559_o = n25544_o;
      4'b0100: n25559_o = n25478_o;
      4'b0010: n25559_o = n25348_o;
      4'b0001: n25559_o = n25232_o;
      default: n25559_o = 1'bX;
    endcase
  assign n25560_o = r1[135];
  assign n25561_o = n25085_o[133];
  assign n25562_o = r1[135];
  /* dcache.vhdl:1373:21  */
  assign n25563_o = n25084_o ? n25561_o : n25562_o;
  /* dcache.vhdl:1346:17  */
  assign n25564_o = n25044_o ? n25560_o : n25563_o;
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25566_o = n25564_o;
      4'b0100: n25566_o = n25564_o;
      4'b0010: n25566_o = n25564_o;
      4'b0001: n25566_o = 1'b1;
      default: n25566_o = 1'bX;
    endcase
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25568_o = n25546_o;
      4'b0100: n25568_o = n25513_o;
      4'b0010: n25568_o = n25381_o;
      4'b0001: n25568_o = n25235_o;
      default: n25568_o = 2'bX;
    endcase
  assign n25569_o = r1[336];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25571_o = n25569_o;
      4'b0100: n25571_o = n25569_o;
      4'b0010: n25571_o = n25569_o;
      4'b0001: n25571_o = n25107_o;
      default: n25571_o = 1'bX;
    endcase
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25573_o = 1'b0;
      4'b0100: n25573_o = n25472_o;
      4'b0010: n25573_o = 1'b0;
      4'b0001: n25573_o = n25237_o;
      default: n25573_o = 1'bX;
    endcase
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25575_o = n25043_o;
      4'b0100: n25575_o = n25043_o;
      4'b0010: n25575_o = n25043_o;
      4'b0001: n25575_o = n25239_o;
      default: n25575_o = 1'bX;
    endcase
  assign n25576_o = n25494_o[0];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25578_o = n25547_o;
      4'b0100: n25578_o = n25576_o;
      4'b0010: n25578_o = n25349_o;
      4'b0001: n25578_o = n25241_o;
      default: n25578_o = 1'bX;
    endcase
  assign n25579_o = n25104_o[4:0];
  assign n25580_o = n25299_o[4:0];
  assign n25581_o = n25494_o[5:1];
  assign n25582_o = r1[344:340];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25584_o = n25582_o;
      4'b0100: n25584_o = n25581_o;
      4'b0010: n25584_o = n25580_o;
      4'b0001: n25584_o = n25579_o;
      default: n25584_o = 5'bX;
    endcase
  assign n25585_o = n25104_o[28:5];
  assign n25586_o = n25299_o[28:5];
  assign n25587_o = r1[368:345];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25589_o = n25587_o;
      4'b0100: n25589_o = n25587_o;
      4'b0010: n25589_o = n25586_o;
      4'b0001: n25589_o = n25585_o;
      default: n25589_o = 24'bX;
    endcase
  assign n25590_o = n25443_o[63:0];
  assign n25591_o = r1[432:369];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25593_o = n25591_o;
      4'b0100: n25593_o = n25590_o;
      4'b0010: n25593_o = n25591_o;
      4'b0001: n25593_o = n25106_o;
      default: n25593_o = 64'bX;
    endcase
  assign n25594_o = n25443_o[71:64];
  assign n25595_o = r1[440:433];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25597_o = n25595_o;
      4'b0100: n25597_o = n25594_o;
      4'b0010: n25597_o = n25595_o;
      4'b0001: n25597_o = n25105_o;
      default: n25597_o = 8'bX;
    endcase
  assign n25598_o = n25522_o[0];
  assign n25599_o = n25550_o[0];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25601_o = n25599_o;
      4'b0100: n25601_o = n25598_o;
      4'b0010: n25601_o = n25383_o;
      4'b0001: n25601_o = n25244_o;
      default: n25601_o = 1'bX;
    endcase
  assign n25602_o = n25522_o[1];
  assign n25603_o = n25550_o[1];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25605_o = n25603_o;
      4'b0100: n25605_o = n25602_o;
      4'b0010: n25605_o = n25281_o;
      4'b0001: n25605_o = n25247_o;
      default: n25605_o = 1'bX;
    endcase
  assign n25606_o = r1[443];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25608_o = n25606_o;
      4'b0100: n25608_o = n25606_o;
      4'b0010: n25608_o = n25606_o;
      4'b0001: n25608_o = n25250_o;
      default: n25608_o = 1'bX;
    endcase
  assign n25609_o = r1[491:444];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25611_o = n25609_o;
      4'b0100: n25611_o = n25609_o;
      4'b0010: n25611_o = n25609_o;
      4'b0001: n25611_o = n25149_o;
      default: n25611_o = 48'bX;
    endcase
  assign n25612_o = r1[496:492];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25614_o = n25612_o;
      4'b0100: n25614_o = n25483_o;
      4'b0010: n25614_o = n25411_o;
      4'b0001: n25614_o = n25122_o;
      default: n25614_o = 5'bX;
    endcase
  assign n25615_o = r1[498:497];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25617_o = n25615_o;
      4'b0100: n25617_o = n25615_o;
      4'b0010: n25617_o = n25615_o;
      4'b0001: n25617_o = n25114_o;
      default: n25617_o = 2'bX;
    endcase
  assign n25618_o = r1[501:499];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25620_o = n25618_o;
      4'b0100: n25620_o = n25618_o;
      4'b0010: n25620_o = n25618_o;
      4'b0001: n25620_o = n25142_o;
      default: n25620_o = 3'bX;
    endcase
  assign n25621_o = n25413_o[0];
  assign n25622_o = r1[502];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25624_o = n25622_o;
      4'b0100: n25624_o = n25622_o;
      4'b0010: n25624_o = n25621_o;
      4'b0001: n25624_o = 1'b0;
      default: n25624_o = 1'bX;
    endcase
  assign n25625_o = n25413_o[1];
  assign n25626_o = r1[503];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25628_o = n25626_o;
      4'b0100: n25628_o = n25626_o;
      4'b0010: n25628_o = n25625_o;
      4'b0001: n25628_o = 1'b0;
      default: n25628_o = 1'bX;
    endcase
  assign n25629_o = n25413_o[2];
  assign n25630_o = r1[504];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25632_o = n25630_o;
      4'b0100: n25632_o = n25630_o;
      4'b0010: n25632_o = n25629_o;
      4'b0001: n25632_o = 1'b0;
      default: n25632_o = 1'bX;
    endcase
  assign n25633_o = n25413_o[3];
  assign n25634_o = r1[505];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25636_o = n25634_o;
      4'b0100: n25636_o = n25634_o;
      4'b0010: n25636_o = n25633_o;
      4'b0001: n25636_o = 1'b0;
      default: n25636_o = 1'bX;
    endcase
  assign n25637_o = n25413_o[4];
  assign n25638_o = r1[506];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25640_o = n25638_o;
      4'b0100: n25640_o = n25638_o;
      4'b0010: n25640_o = n25637_o;
      4'b0001: n25640_o = 1'b0;
      default: n25640_o = 1'bX;
    endcase
  assign n25641_o = n25413_o[5];
  assign n25642_o = r1[507];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25644_o = n25642_o;
      4'b0100: n25644_o = n25642_o;
      4'b0010: n25644_o = n25641_o;
      4'b0001: n25644_o = 1'b0;
      default: n25644_o = 1'bX;
    endcase
  assign n25645_o = n25413_o[6];
  assign n25646_o = r1[508];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25648_o = n25646_o;
      4'b0100: n25648_o = n25646_o;
      4'b0010: n25648_o = n25645_o;
      4'b0001: n25648_o = 1'b0;
      default: n25648_o = 1'bX;
    endcase
  assign n25649_o = n25413_o[7];
  assign n25650_o = r1[509];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25652_o = n25650_o;
      4'b0100: n25652_o = n25650_o;
      4'b0010: n25652_o = n25649_o;
      4'b0001: n25652_o = 1'b0;
      default: n25652_o = 1'bX;
    endcase
  assign n25653_o = r1[512:510];
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25655_o = n25653_o;
      4'b0100: n25655_o = n25432_o;
      4'b0010: n25655_o = n25653_o;
      4'b0001: n25655_o = n25253_o;
      default: n25655_o = 3'bX;
    endcase
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25657_o = 1'b0;
      4'b0100: n25657_o = n25484_o;
      4'b0010: n25657_o = 1'b0;
      4'b0001: n25657_o = 1'b0;
      default: n25657_o = 1'bX;
    endcase
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25659_o = 1'b0;
      4'b0100: n25659_o = n25523_o;
      4'b0010: n25659_o = 1'b0;
      4'b0001: n25659_o = 1'b0;
      default: n25659_o = 1'bX;
    endcase
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25661_o = n25539_o;
      4'b0100: n25661_o = n25485_o;
      4'b0010: n25661_o = n25346_o;
      4'b0001: n25661_o = n25255_o;
      default: n25661_o = 1'bX;
    endcase
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25663_o = n25552_o;
      4'b0100: n25663_o = n25018_o;
      4'b0010: n25663_o = n25351_o;
      4'b0001: n25663_o = n25257_o;
      default: n25663_o = 1'bX;
    endcase
  assign n25664_o = r1[136];
  assign n25665_o = n25085_o[134];
  assign n25666_o = r1[136];
  /* dcache.vhdl:1373:21  */
  assign n25667_o = n25084_o ? n25665_o : n25666_o;
  /* dcache.vhdl:1346:17  */
  assign n25668_o = n25044_o ? n25664_o : n25667_o;
  assign n25669_o = r1[134:2];
  assign n25670_o = n25085_o[132:0];
  assign n25671_o = r1[134:2];
  /* dcache.vhdl:1373:21  */
  assign n25672_o = n25084_o ? n25670_o : n25671_o;
  /* dcache.vhdl:1346:17  */
  assign n25673_o = n25044_o ? n25669_o : n25672_o;
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25675_o = 1'b0;
      4'b0100: n25675_o = 1'b0;
      4'b0010: n25675_o = 1'b0;
      4'b0001: n25675_o = n25259_o;
      default: n25675_o = 1'bX;
    endcase
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25677_o = 1'b0;
      4'b0100: n25677_o = 1'b0;
      4'b0010: n25677_o = 1'b0;
      4'b0001: n25677_o = n25261_o;
      default: n25677_o = 1'bX;
    endcase
  /* dcache.vhdl:1381:17  */
  always @*
    case (n25555_o)
      4'b1000: n25679_o = 1'b0;
      4'b0100: n25679_o = 1'b0;
      4'b0010: n25679_o = n25384_o;
      4'b0001: n25679_o = 1'b0;
      default: n25679_o = 1'bX;
    endcase
  assign n25685_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* dcache.vhdl:1293:13  */
  assign n25686_o = rst ? n25685_o : n25557_o;
  assign n25687_o = {n25668_o, n25566_o, n25673_o};
  assign n25688_o = {n25661_o, n25659_o, n25657_o, n25655_o, n25652_o, n25648_o, n25644_o, n25640_o, n25636_o, n25632_o, n25628_o, n25624_o, n25620_o, n25617_o, n25614_o, n25611_o, n25608_o, n25605_o, n25601_o, n25597_o, n25593_o, n25589_o, n25584_o, n25578_o, n25575_o, n25573_o, n25571_o, n25568_o};
  assign n25689_o = {29'b00000000000000000000000000000, 1'b0};
  assign n25690_o = {1'b0, 1'b0};
  /* dcache.vhdl:1293:13  */
  assign n25691_o = rst ? 1'b0 : n25559_o;
  assign n25692_o = r1[136:2];
  /* dcache.vhdl:1293:13  */
  assign n25693_o = rst ? n25692_o : n25687_o;
  assign n25694_o = n25688_o[1:0];
  /* dcache.vhdl:1293:13  */
  assign n25695_o = rst ? 2'b00 : n25694_o;
  assign n25696_o = n25688_o[4:2];
  assign n25697_o = r1[338:336];
  /* dcache.vhdl:1293:13  */
  assign n25698_o = rst ? n25697_o : n25696_o;
  assign n25699_o = n25688_o[34:5];
  /* dcache.vhdl:1293:13  */
  assign n25700_o = rst ? n25689_o : n25699_o;
  assign n25701_o = n25688_o[106:35];
  assign n25702_o = r1[440:369];
  /* dcache.vhdl:1293:13  */
  assign n25703_o = rst ? n25702_o : n25701_o;
  assign n25704_o = n25688_o[108:107];
  /* dcache.vhdl:1293:13  */
  assign n25705_o = rst ? n25690_o : n25704_o;
  assign n25706_o = n25688_o[180:109];
  assign n25707_o = r1[514:443];
  /* dcache.vhdl:1293:13  */
  assign n25708_o = rst ? n25707_o : n25706_o;
  assign n25709_o = n25688_o[181];
  /* dcache.vhdl:1293:13  */
  assign n25710_o = rst ? 1'b0 : n25709_o;
  /* dcache.vhdl:1293:13  */
  assign n25711_o = rst ? 1'b0 : n25663_o;
  assign n25712_o = {n25679_o, n25677_o, n25675_o};
  assign n25713_o = {1'b0, 1'b0, 1'b0};
  /* dcache.vhdl:1293:13  */
  assign n25714_o = rst ? n25713_o : n25712_o;
  assign n25720_o = {n25710_o, n25708_o, n25705_o, n25703_o, n25700_o, n25698_o, n25695_o};
  assign n25729_o = {tlb_miss, n25714_o};
  /* dcache.vhdl:1293:13  */
  assign n25739_o = ~rst;
  /* dcache.vhdl:1293:13  */
  assign n25740_o = n25739_o & n25032_o;
  /* dcache.vhdl:1286:9  */
  always @(posedge clk)
    n25744_q <= n25686_o;
  /* dcache.vhdl:719:9  */
  always @(posedge clk)
    n25745_q <= n24103_o;
  /* dcache.vhdl:723:13  */
  assign n25746_o = ~n24025_o;
  /* dcache.vhdl:728:13  */
  assign n25747_o = ~n24020_o;
  /* dcache.vhdl:723:13  */
  assign n25748_o = n25746_o & n25747_o;
  /* dcache.vhdl:723:13  */
  assign n25749_o = n25748_o & n24022_o;
  /* dcache.vhdl:723:13  */
  assign n25752_o = ~n24025_o;
  /* dcache.vhdl:728:13  */
  assign n25753_o = ~n24020_o;
  /* dcache.vhdl:723:13  */
  assign n25754_o = n25752_o & n25753_o;
  /* dcache.vhdl:723:13  */
  assign n25755_o = n25754_o & n24022_o;
  /* dcache.vhdl:561:9  */
  always @(posedge clk)
    n25758_q <= n23835_o;
  /* dcache.vhdl:561:9  */
  always @(posedge clk)
    n25759_q <= n23837_o;
  /* dcache.vhdl:1286:9  */
  always @(posedge clk)
    n25760_q <= n25711_o;
  /* dcache.vhdl:1286:9  */
  always @(posedge clk)
    n25761_q <= n25720_o;
  /* dcache.vhdl:1286:9  */
  always @(posedge clk)
    n25762_q <= n25693_o;
  /* dcache.vhdl:1286:9  */
  always @(posedge clk)
    n25763_q <= n25691_o;
  /* dcache.vhdl:1181:9  */
  always @(posedge clk)
    n25764_q <= n24962_o;
  /* dcache.vhdl:1181:9  */
  always @(posedge clk)
    n25765_q <= n24954_o;
  /* dcache.vhdl:1181:9  */
  always @(posedge clk)
    n25766_q <= n24961_o;
  /* dcache.vhdl:1181:9  */
  assign n25767_o = r1[1];
  /* dcache.vhdl:1181:9  */
  assign n25768_o = r0_valid ? n24701_o : n25767_o;
  /* dcache.vhdl:1181:9  */
  always @(posedge clk)
    n25769_q <= n25768_o;
  /* dcache.vhdl:1181:9  */
  assign n25770_o = {n25764_q, n25760_q, n25765_q, n25761_q, n25766_q, n25762_q, n25769_q, n25763_q};
  /* dcache.vhdl:1286:9  */
  always @(posedge clk)
    n25771_q <= n25729_o;
  /* dcache.vhdl:719:9  */
  always @(posedge clk)
    n25772_q <= n24022_o;
  /* dcache.vhdl:719:9  */
  assign n25773_o = {n25772_q, n25771_q};
  /* dcache.vhdl:1021:9  */
  always @(posedge clk)
    n25774_q <= n24635_o;
  /* dcache.vhdl:621:9  */
  assign n25783_o = n23864_o ? n25805_o : tlb_valid_way;
  /* dcache.vhdl:621:9  */
  always @(posedge clk)
    n25784_q <= n25783_o;
  /* dcache.vhdl:621:9  */
  assign n25785_o = {maybe_tlb_plrus_tlb_plrus_n1_tlb_plru_out, maybe_tlb_plrus_tlb_plrus_n2_tlb_plru_out};
  /* dcache.vhdl:806:9  */
  always @(posedge clk)
    n25787_q <= n24211_o;
  /* dcache.vhdl:806:9  */
  always @(posedge clk)
    n25788_q <= n24191_o;
  /* dcache.vhdl:806:9  */
  always @(posedge clk)
    n25789_q <= n24197_o;
  /* dcache.vhdl:806:9  */
  assign n25790_o = {n24644_o, n24643_o, n24642_o, n24640_o, n24639_o};
  assign n25791_o = {n24647_o, n24646_o, n24645_o, 1'b0};
  /* dcache.vhdl:632:42  */
  reg [101:0] dtlb_tags[1:0] ; // memory
  always @(posedge clk)
    if (n23864_o)
      n25794_data <= dtlb_tags[n23862_o];
  always @(posedge clk)
    if (n25749_o)
      dtlb_tags[tlb_req_index] <= n25836_o;
  /* dcache.vhdl:621:9  */
  /* dcache.vhdl:741:27  */
  /* dcache.vhdl:633:42  */
  reg [127:0] dtlb_ptes[1:0] ; // memory
  always @(posedge clk)
    if (n23864_o)
      n25796_data <= dtlb_ptes[n23862_o];
  always @(posedge clk)
    if (n25755_o)
      dtlb_ptes[tlb_req_index] <= n25843_o;
  /* dcache.vhdl:621:9  */
  /* dcache.vhdl:744:27  */
  /* dcache.vhdl:798:41  */
  reg [47:0] cache_tags[3:0] ; // memory
  always @(posedge clk)
    if (1'b1)
      n25799_data <= cache_tags[n24180_o];
  always @(posedge clk)
    if (1'b1)
      n25801_data <= cache_tags[n24147_o];
  always @(posedge clk)
    if (n25740_o)
      cache_tags[n25033_o] <= n25037_o;
  /* dcache.vhdl:798:41  */
  /* dcache.vhdl:808:40  */
  /* dcache.vhdl:1336:43  */
  /* dcache.vhdl:723:13  */
  assign n25803_o = dtlb_valids[1:0];
  /* dcache.vhdl:723:13  */
  assign n25804_o = dtlb_valids[3:2];
  /* dcache.vhdl:631:45  */
  assign n25805_o = n23866_o ? n25804_o : n25803_o;
  /* dcache.vhdl:631:45  */
  assign n25806_o = tlb_pte_way[63:0];
  /* dcache.vhdl:631:46  */
  assign n25807_o = tlb_pte_way[127:64];
  /* dcache.vhdl:528:20  */
  assign n25808_o = n23945_o ? n25807_o : n25806_o;
  /* dcache.vhdl:730:47  */
  assign n25809_o = {n24029_o, tlb_hit_way};
  /* dcache.vhdl:730:21  */
  assign n25810_o = n25809_o[1];
  /* dcache.vhdl:730:21  */
  assign n25811_o = ~n25810_o;
  /* dcache.vhdl:730:21  */
  assign n25812_o = n25809_o[0];
  /* dcache.vhdl:730:21  */
  assign n25813_o = ~n25812_o;
  /* dcache.vhdl:730:21  */
  assign n25814_o = n25811_o & n25813_o;
  /* dcache.vhdl:730:21  */
  assign n25815_o = n25811_o & n25812_o;
  /* dcache.vhdl:730:21  */
  assign n25816_o = n25810_o & n25813_o;
  /* dcache.vhdl:730:21  */
  assign n25817_o = n25810_o & n25812_o;
  /* dcache.vhdl:1336:43  */
  assign n25818_o = dtlb_valids[0];
  /* dcache.vhdl:730:21  */
  assign n25819_o = n25814_o ? 1'b0 : n25818_o;
  /* dcache.vhdl:153:12  */
  assign n25820_o = dtlb_valids[1];
  /* dcache.vhdl:730:21  */
  assign n25821_o = n25815_o ? 1'b0 : n25820_o;
  /* dcache.vhdl:633:41  */
  assign n25822_o = dtlb_valids[2];
  /* dcache.vhdl:730:21  */
  assign n25823_o = n25816_o ? 1'b0 : n25822_o;
  /* dcache.vhdl:633:42  */
  assign n25824_o = dtlb_valids[3];
  /* dcache.vhdl:730:21  */
  assign n25825_o = n25817_o ? 1'b0 : n25824_o;
  /* dcache.vhdl:744:27  */
  assign n25826_o = {n25825_o, n25823_o, n25821_o, n25819_o};
  /* dcache.vhdl:730:48  */
  assign n25827_o = tlb_plru_victim[0];
  /* dcache.vhdl:730:33  */
  assign n25828_o = tlb_plru_victim[1];
  /* dcache.vhdl:736:68  */
  assign n25829_o = n24037_o ? n25828_o : n25827_o;
  /* dcache.vhdl:520:9  */
  assign n25830_o = n24041_o;
  /* dcache.vhdl:520:9  */
  assign n25831_o = ~n25830_o;
  /* dcache.vhdl:744:27  */
  assign n25832_o = tlb_tag_way[50:0];
  /* dcache.vhdl:520:9  */
  assign n25833_o = n25831_o ? n24042_o : n25832_o;
  /* dcache.vhdl:741:17  */
  assign n25834_o = tlb_tag_way[101:51];
  /* dcache.vhdl:520:9  */
  assign n25835_o = n25830_o ? n24042_o : n25834_o;
  /* dcache.vhdl:621:9  */
  assign n25836_o = {n25835_o, n25833_o};
  /* dcache.vhdl:535:9  */
  assign n25837_o = n24041_o;
  /* dcache.vhdl:535:9  */
  assign n25838_o = ~n25837_o;
  /* dcache.vhdl:632:42  */
  assign n25839_o = tlb_pte_way[63:0];
  /* dcache.vhdl:535:9  */
  assign n25840_o = n25838_o ? n24063_o : n25839_o;
  /* dcache.vhdl:741:27  */
  assign n25841_o = tlb_pte_way[127:64];
  /* dcache.vhdl:535:9  */
  assign n25842_o = n25837_o ? n24063_o : n25841_o;
  /* dcache.vhdl:1141:28  */
  assign n25843_o = {n25842_o, n25840_o};
  /* dcache.vhdl:745:43  */
  assign n25844_o = {n24082_o, n24041_o};
  /* dcache.vhdl:745:17  */
  assign n25845_o = n25844_o[1];
  /* dcache.vhdl:745:17  */
  assign n25846_o = ~n25845_o;
  /* dcache.vhdl:745:17  */
  assign n25847_o = n25844_o[0];
  /* dcache.vhdl:745:17  */
  assign n25848_o = ~n25847_o;
  /* dcache.vhdl:745:17  */
  assign n25849_o = n25846_o & n25848_o;
  /* dcache.vhdl:745:17  */
  assign n25850_o = n25846_o & n25847_o;
  /* dcache.vhdl:745:17  */
  assign n25851_o = n25845_o & n25848_o;
  /* dcache.vhdl:745:17  */
  assign n25852_o = n25845_o & n25847_o;
  /* dcache.vhdl:49:9  */
  assign n25853_o = dtlb_valids[0];
  /* dcache.vhdl:745:17  */
  assign n25854_o = n25849_o ? 1'b1 : n25853_o;
  /* dcache.vhdl:44:9  */
  assign n25855_o = dtlb_valids[1];
  /* dcache.vhdl:745:17  */
  assign n25856_o = n25850_o ? 1'b1 : n25855_o;
  /* dcache.vhdl:37:9  */
  assign n25857_o = dtlb_valids[2];
  /* dcache.vhdl:745:17  */
  assign n25858_o = n25851_o ? 1'b1 : n25857_o;
  assign n25859_o = dtlb_valids[3];
  /* dcache.vhdl:745:17  */
  assign n25860_o = n25852_o ? 1'b1 : n25859_o;
  assign n25861_o = {n25860_o, n25858_o, n25856_o, n25854_o};
  /* dcache.vhdl:745:44  */
  assign n25862_o = cache_valids[0];
  /* dcache.vhdl:745:29  */
  assign n25863_o = cache_valids[1];
  /* dcache.vhdl:745:17  */
  assign n25864_o = cache_valids[2];
  /* dcache.vhdl:1021:9  */
  assign n25865_o = cache_valids[3];
  /* dcache.vhdl:864:60  */
  assign n25866_o = n24287_o[1:0];
  /* dcache.vhdl:864:60  */
  always @*
    case (n25866_o)
      2'b00: n25867_o = n25862_o;
      2'b01: n25867_o = n25863_o;
      2'b10: n25867_o = n25864_o;
      2'b11: n25867_o = n25865_o;
    endcase
  /* dcache.vhdl:864:60  */
  assign n25868_o = cache_valids[0];
  /* dcache.vhdl:864:50  */
  assign n25869_o = cache_valids[1];
  /* dcache.vhdl:1286:9  */
  assign n25870_o = cache_valids[2];
  assign n25871_o = cache_valids[3];
  /* dcache.vhdl:864:60  */
  assign n25872_o = n24335_o[1:0];
  /* dcache.vhdl:864:60  */
  always @*
    case (n25872_o)
      2'b00: n25873_o = n25868_o;
      2'b01: n25873_o = n25869_o;
      2'b10: n25873_o = n25870_o;
      2'b11: n25873_o = n25871_o;
    endcase
  /* dcache.vhdl:864:60  */
  assign n25874_o = n24361_o[0];
  /* dcache.vhdl:864:50  */
  assign n25875_o = n24361_o[1];
  /* dcache.vhdl:880:34  */
  assign n25876_o = tlb_hit_way ? n25875_o : n25874_o;
  /* dcache.vhdl:880:34  */
  assign n25877_o = n24367_o[0];
  /* dcache.vhdl:880:35  */
  assign n25878_o = n24367_o[1];
  /* dcache.vhdl:882:41  */
  assign n25879_o = tlb_hit_way ? n25878_o : n25877_o;
  /* dcache.vhdl:882:41  */
  assign n25880_o = n24370_o[0];
  /* dcache.vhdl:882:42  */
  assign n25881_o = n24370_o[1];
  /* dcache.vhdl:883:41  */
  assign n25882_o = tlb_hit_way ? n25881_o : n25880_o;
  /* dcache.vhdl:883:41  */
  assign n25883_o = cache_valids[0];
  /* dcache.vhdl:883:42  */
  assign n25884_o = cache_valids[1];
  /* dcache.vhdl:1293:13  */
  assign n25885_o = cache_valids[2];
  /* dcache.vhdl:1293:13  */
  assign n25886_o = cache_valids[3];
  /* dcache.vhdl:888:56  */
  assign n25887_o = n24387_o[1:0];
  /* dcache.vhdl:888:56  */
  always @*
    case (n25887_o)
      2'b00: n25888_o = n25883_o;
      2'b01: n25888_o = n25884_o;
      2'b10: n25888_o = n25885_o;
      2'b11: n25888_o = n25886_o;
    endcase
  /* dcache.vhdl:888:56  */
  assign n25889_o = r1[502];
  /* dcache.vhdl:888:46  */
  assign n25890_o = r1[503];
  assign n25891_o = r1[504];
  /* dcache.vhdl:1381:17  */
  assign n25892_o = r1[505];
  assign n25893_o = r1[506];
  assign n25894_o = r1[507];
  assign n25895_o = r1[508];
  assign n25896_o = r1[509];
  /* dcache.vhdl:935:55  */
  assign n25897_o = n24479_o[1:0];
  /* dcache.vhdl:935:55  */
  always @*
    case (n25897_o)
      2'b00: n25898_o = n25889_o;
      2'b01: n25898_o = n25890_o;
      2'b10: n25898_o = n25891_o;
      2'b11: n25898_o = n25892_o;
    endcase
  /* dcache.vhdl:935:55  */
  assign n25899_o = n24479_o[1:0];
  /* dcache.vhdl:935:55  */
  always @*
    case (n25899_o)
      2'b00: n25900_o = n25893_o;
      2'b01: n25900_o = n25894_o;
      2'b10: n25900_o = n25895_o;
      2'b11: n25900_o = n25896_o;
    endcase
  /* dcache.vhdl:935:55  */
  assign n25901_o = n24479_o[2];
  /* dcache.vhdl:935:55  */
  assign n25902_o = n25901_o ? n25900_o : n25898_o;
  /* dcache.vhdl:1328:25  */
  assign n25903_o = n25027_o[1];
  /* dcache.vhdl:1328:25  */
  assign n25904_o = ~n25903_o;
  /* dcache.vhdl:1328:25  */
  assign n25905_o = n25027_o[0];
  /* dcache.vhdl:1328:25  */
  assign n25906_o = ~n25905_o;
  /* dcache.vhdl:1328:25  */
  assign n25907_o = n25904_o & n25906_o;
  /* dcache.vhdl:1328:25  */
  assign n25908_o = n25904_o & n25905_o;
  /* dcache.vhdl:1328:25  */
  assign n25909_o = n25903_o & n25906_o;
  /* dcache.vhdl:1328:25  */
  assign n25910_o = n25903_o & n25905_o;
  assign n25911_o = cache_valids[0];
  /* dcache.vhdl:1328:25  */
  assign n25912_o = n25907_o ? 1'b0 : n25911_o;
  assign n25913_o = cache_valids[1];
  /* dcache.vhdl:1328:25  */
  assign n25914_o = n25908_o ? 1'b0 : n25913_o;
  assign n25915_o = cache_valids[2];
  /* dcache.vhdl:1328:25  */
  assign n25916_o = n25909_o ? 1'b0 : n25915_o;
  /* dcache.vhdl:483:14  */
  assign n25917_o = cache_valids[3];
  /* dcache.vhdl:1328:25  */
  assign n25918_o = n25910_o ? 1'b0 : n25917_o;
  /* dcache.vhdl:483:14  */
  assign n25919_o = {n25918_o, n25916_o, n25914_o, n25912_o};
  /* dcache.vhdl:1481:25  */
  assign n25920_o = n25308_o[2];
  /* dcache.vhdl:1481:25  */
  assign n25921_o = ~n25920_o;
  /* dcache.vhdl:1481:25  */
  assign n25922_o = n25308_o[1];
  /* dcache.vhdl:1481:25  */
  assign n25923_o = ~n25922_o;
  /* dcache.vhdl:1481:25  */
  assign n25924_o = n25921_o & n25923_o;
  /* dcache.vhdl:1481:25  */
  assign n25925_o = n25921_o & n25922_o;
  /* dcache.vhdl:1481:25  */
  assign n25926_o = n25920_o & n25923_o;
  /* dcache.vhdl:1481:25  */
  assign n25927_o = n25920_o & n25922_o;
  /* dcache.vhdl:1481:25  */
  assign n25928_o = n25308_o[0];
  /* dcache.vhdl:1481:25  */
  assign n25929_o = ~n25928_o;
  /* dcache.vhdl:1481:25  */
  assign n25930_o = n25924_o & n25929_o;
  /* dcache.vhdl:1481:25  */
  assign n25931_o = n25924_o & n25928_o;
  /* dcache.vhdl:1481:25  */
  assign n25932_o = n25925_o & n25929_o;
  /* dcache.vhdl:1481:25  */
  assign n25933_o = n25925_o & n25928_o;
  /* dcache.vhdl:1481:25  */
  assign n25934_o = n25926_o & n25929_o;
  /* dcache.vhdl:1481:25  */
  assign n25935_o = n25926_o & n25928_o;
  /* dcache.vhdl:1481:25  */
  assign n25936_o = n25927_o & n25929_o;
  /* dcache.vhdl:1481:25  */
  assign n25937_o = n25927_o & n25928_o;
  /* dcache.vhdl:441:14  */
  assign n25938_o = n25310_o[0];
  /* dcache.vhdl:1481:25  */
  assign n25939_o = n25930_o ? 1'b1 : n25938_o;
  assign n25940_o = n25310_o[1];
  /* dcache.vhdl:1481:25  */
  assign n25941_o = n25931_o ? 1'b1 : n25940_o;
  assign n25942_o = n25310_o[2];
  /* dcache.vhdl:1481:25  */
  assign n25943_o = n25932_o ? 1'b1 : n25942_o;
  assign n25944_o = n25310_o[3];
  /* dcache.vhdl:1481:25  */
  assign n25945_o = n25933_o ? 1'b1 : n25944_o;
  assign n25946_o = n25310_o[4];
  /* dcache.vhdl:1481:25  */
  assign n25947_o = n25934_o ? 1'b1 : n25946_o;
  /* dcache.vhdl:467:14  */
  assign n25948_o = n25310_o[5];
  /* dcache.vhdl:1481:25  */
  assign n25949_o = n25935_o ? 1'b1 : n25948_o;
  /* dcache.vhdl:467:14  */
  assign n25950_o = n25310_o[6];
  /* dcache.vhdl:1481:25  */
  assign n25951_o = n25936_o ? 1'b1 : n25950_o;
  /* dcache.vhdl:455:14  */
  assign n25952_o = n25310_o[7];
  /* dcache.vhdl:1481:25  */
  assign n25953_o = n25937_o ? 1'b1 : n25952_o;
  /* dcache.vhdl:455:14  */
  assign n25954_o = {n25953_o, n25951_o, n25949_o, n25947_o, n25945_o, n25943_o, n25941_o, n25939_o};
  /* dcache.vhdl:1506:29  */
  assign n25955_o = n25372_o[1];
  /* dcache.vhdl:1506:29  */
  assign n25956_o = ~n25955_o;
  /* dcache.vhdl:1506:29  */
  assign n25957_o = n25372_o[0];
  /* dcache.vhdl:1506:29  */
  assign n25958_o = ~n25957_o;
  /* dcache.vhdl:1506:29  */
  assign n25959_o = n25956_o & n25958_o;
  /* dcache.vhdl:1506:29  */
  assign n25960_o = n25956_o & n25957_o;
  /* dcache.vhdl:1506:29  */
  assign n25961_o = n25955_o & n25958_o;
  /* dcache.vhdl:1506:29  */
  assign n25962_o = n25955_o & n25957_o;
  /* dcache.vhdl:495:14  */
  assign n25963_o = n25031_o[0];
  /* dcache.vhdl:1506:29  */
  assign n25964_o = n25959_o ? 1'b1 : n25963_o;
  /* dcache.vhdl:450:30  */
  assign n25965_o = n25031_o[1];
  /* dcache.vhdl:1506:29  */
  assign n25966_o = n25960_o ? 1'b1 : n25965_o;
  assign n25967_o = n25031_o[2];
  /* dcache.vhdl:1506:29  */
  assign n25968_o = n25961_o ? 1'b1 : n25967_o;
  /* dcache.vhdl:447:14  */
  assign n25969_o = n25031_o[3];
  /* dcache.vhdl:1506:29  */
  assign n25970_o = n25962_o ? 1'b1 : n25969_o;
  /* dcache.vhdl:447:14  */
  assign n25971_o = {n25970_o, n25968_o, n25966_o, n25964_o};
endmodule

module mmu
  (input  clk,
   input  rst,
   input  l_in_valid,
   input  l_in_tlbie,
   input  l_in_slbia,
   input  l_in_mtspr,
   input  l_in_iside,
   input  l_in_load,
   input  l_in_priv,
   input  [9:0] l_in_sprn,
   input  [63:0] l_in_addr,
   input  [63:0] l_in_rs,
   input  d_in_stall,
   input  d_in_done,
   input  d_in_err,
   input  [63:0] d_in_data,
   output l_out_done,
   output l_out_err,
   output l_out_invalid,
   output l_out_badtree,
   output l_out_segerr,
   output l_out_perm_error,
   output l_out_rc_error,
   output [63:0] l_out_sprval,
   output d_out_valid,
   output d_out_tlbie,
   output d_out_doall,
   output d_out_tlbld,
   output [63:0] d_out_addr,
   output [63:0] d_out_pte,
   output i_out_tlbld,
   output i_out_tlbie,
   output i_out_doall,
   output [63:0] i_out_addr,
   output [63:0] i_out_pte);
  wire [144:0] n22421_o;
  wire n22423_o;
  wire n22424_o;
  wire n22425_o;
  wire n22426_o;
  wire n22427_o;
  wire n22428_o;
  wire n22429_o;
  wire [63:0] n22430_o;
  wire n22432_o;
  wire n22433_o;
  wire n22434_o;
  wire n22435_o;
  wire [63:0] n22436_o;
  wire [63:0] n22437_o;
  wire [66:0] n22438_o;
  wire n22440_o;
  wire n22441_o;
  wire n22442_o;
  wire [63:0] n22443_o;
  wire [63:0] n22444_o;
  wire [501:0] r;
  wire [501:0] rin;
  wire [15:0] addrsh;
  wire [15:0] mask;
  wire [43:0] finalmask;
  wire [63:0] n22445_o;
  wire n22446_o;
  wire [63:0] n22447_o;
  wire [31:0] n22448_o;
  wire [63:0] n22450_o;
  wire [99:0] n22469_o;
  wire n22470_o;
  wire n22471_o;
  wire [67:0] n22472_o;
  wire [67:0] n22473_o;
  wire [67:0] n22474_o;
  wire [99:0] n22475_o;
  wire [99:0] n22476_o;
  wire [65:0] n22477_o;
  wire [65:0] n22478_o;
  wire [65:0] n22479_o;
  wire n22480_o;
  wire n22481_o;
  wire [63:0] n22482_o;
  wire [63:0] n22483_o;
  wire [63:0] n22484_o;
  wire n22485_o;
  wire n22486_o;
  wire [63:0] n22487_o;
  wire [63:0] n22488_o;
  wire [63:0] n22489_o;
  wire n22490_o;
  wire n22491_o;
  wire [135:0] n22492_o;
  wire [135:0] n22493_o;
  wire [135:0] n22494_o;
  wire [501:0] n22495_o;
  wire [1:0] n22502_o;
  wire [30:0] n22503_o;
  wire n22505_o;
  wire [30:0] n22506_o;
  wire n22508_o;
  wire [17:0] n22509_o;
  wire [30:0] n22511_o;
  wire [1:0] n22512_o;
  reg [30:0] n22513_o;
  wire [1:0] n22514_o;
  wire [18:0] n22515_o;
  wire n22517_o;
  wire [18:0] n22518_o;
  wire n22520_o;
  wire [18:0] n22521_o;
  wire n22523_o;
  wire [18:0] n22524_o;
  wire [2:0] n22525_o;
  reg [18:0] n22526_o;
  wire [1:0] n22527_o;
  wire [15:0] n22528_o;
  wire n22530_o;
  wire [15:0] n22531_o;
  wire n22533_o;
  wire [15:0] n22534_o;
  wire n22536_o;
  wire [15:0] n22537_o;
  wire [2:0] n22538_o;
  reg [15:0] n22539_o;
  wire [4:0] n22543_o;
  wire [30:0] n22544_o;
  wire [31:0] n22545_o;
  wire n22547_o;
  wire n22550_o;
  localparam [15:0] n22551_o = 16'b0000000000011111;
  wire [4:0] n22553_o;
  wire [4:0] n22554_o;
  wire [30:0] n22555_o;
  wire [31:0] n22556_o;
  wire n22558_o;
  wire n22560_o;
  wire n22561_o;
  wire [4:0] n22563_o;
  wire [30:0] n22564_o;
  wire [31:0] n22565_o;
  wire n22567_o;
  wire n22569_o;
  wire n22570_o;
  wire [4:0] n22572_o;
  wire [30:0] n22573_o;
  wire [31:0] n22574_o;
  wire n22576_o;
  wire n22578_o;
  wire n22579_o;
  wire [4:0] n22581_o;
  wire [30:0] n22582_o;
  wire [31:0] n22583_o;
  wire n22585_o;
  wire n22587_o;
  wire n22588_o;
  wire [4:0] n22590_o;
  wire [30:0] n22591_o;
  wire [31:0] n22592_o;
  wire n22594_o;
  wire n22596_o;
  wire n22597_o;
  wire [4:0] n22599_o;
  wire [30:0] n22600_o;
  wire [31:0] n22601_o;
  wire n22603_o;
  wire n22605_o;
  wire n22606_o;
  wire [4:0] n22608_o;
  wire [30:0] n22609_o;
  wire [31:0] n22610_o;
  wire n22612_o;
  wire n22614_o;
  wire n22615_o;
  wire [4:0] n22617_o;
  wire [30:0] n22618_o;
  wire [31:0] n22619_o;
  wire n22621_o;
  wire n22623_o;
  wire n22624_o;
  wire [4:0] n22626_o;
  wire [30:0] n22627_o;
  wire [31:0] n22628_o;
  wire n22630_o;
  wire n22632_o;
  wire n22633_o;
  wire n22634_o;
  wire [4:0] n22635_o;
  wire [30:0] n22636_o;
  wire [31:0] n22637_o;
  wire n22639_o;
  wire n22641_o;
  wire [15:0] n22642_o;
  wire [5:0] n22647_o;
  wire [30:0] n22648_o;
  wire [31:0] n22649_o;
  wire n22651_o;
  wire n22654_o;
  localparam [43:0] n22655_o = 44'b00000000000000000000000000000000000000000000;
  wire [5:0] n22657_o;
  wire [30:0] n22658_o;
  wire [31:0] n22659_o;
  wire n22661_o;
  wire n22663_o;
  wire n22664_o;
  wire [5:0] n22666_o;
  wire [30:0] n22667_o;
  wire [31:0] n22668_o;
  wire n22670_o;
  wire n22672_o;
  wire n22673_o;
  wire [5:0] n22675_o;
  wire [30:0] n22676_o;
  wire [31:0] n22677_o;
  wire n22679_o;
  wire n22681_o;
  wire n22682_o;
  wire [5:0] n22684_o;
  wire [30:0] n22685_o;
  wire [31:0] n22686_o;
  wire n22688_o;
  wire n22690_o;
  wire n22691_o;
  wire [5:0] n22693_o;
  wire [30:0] n22694_o;
  wire [31:0] n22695_o;
  wire n22697_o;
  wire n22699_o;
  wire n22700_o;
  wire [5:0] n22702_o;
  wire [30:0] n22703_o;
  wire [31:0] n22704_o;
  wire n22706_o;
  wire n22708_o;
  wire n22709_o;
  wire [5:0] n22711_o;
  wire [30:0] n22712_o;
  wire [31:0] n22713_o;
  wire n22715_o;
  wire n22717_o;
  wire n22718_o;
  wire [5:0] n22720_o;
  wire [30:0] n22721_o;
  wire [31:0] n22722_o;
  wire n22724_o;
  wire n22726_o;
  wire n22727_o;
  wire [5:0] n22729_o;
  wire [30:0] n22730_o;
  wire [31:0] n22731_o;
  wire n22733_o;
  wire n22735_o;
  wire n22736_o;
  wire [5:0] n22738_o;
  wire [30:0] n22739_o;
  wire [31:0] n22740_o;
  wire n22742_o;
  wire n22744_o;
  wire n22745_o;
  wire [5:0] n22747_o;
  wire [30:0] n22748_o;
  wire [31:0] n22749_o;
  wire n22751_o;
  wire n22753_o;
  wire n22754_o;
  wire [5:0] n22756_o;
  wire [30:0] n22757_o;
  wire [31:0] n22758_o;
  wire n22760_o;
  wire n22762_o;
  wire n22763_o;
  wire [5:0] n22765_o;
  wire [30:0] n22766_o;
  wire [31:0] n22767_o;
  wire n22769_o;
  wire n22771_o;
  wire n22772_o;
  wire [5:0] n22774_o;
  wire [30:0] n22775_o;
  wire [31:0] n22776_o;
  wire n22778_o;
  wire n22780_o;
  wire n22781_o;
  wire [5:0] n22783_o;
  wire [30:0] n22784_o;
  wire [31:0] n22785_o;
  wire n22787_o;
  wire n22789_o;
  wire n22790_o;
  wire [5:0] n22792_o;
  wire [30:0] n22793_o;
  wire [31:0] n22794_o;
  wire n22796_o;
  wire n22798_o;
  wire n22799_o;
  wire [5:0] n22801_o;
  wire [30:0] n22802_o;
  wire [31:0] n22803_o;
  wire n22805_o;
  wire n22807_o;
  wire n22808_o;
  wire [5:0] n22810_o;
  wire [30:0] n22811_o;
  wire [31:0] n22812_o;
  wire n22814_o;
  wire n22816_o;
  wire n22817_o;
  wire [5:0] n22819_o;
  wire [30:0] n22820_o;
  wire [31:0] n22821_o;
  wire n22823_o;
  wire n22825_o;
  wire n22826_o;
  wire [5:0] n22828_o;
  wire [30:0] n22829_o;
  wire [31:0] n22830_o;
  wire n22832_o;
  wire n22834_o;
  wire n22835_o;
  wire [5:0] n22837_o;
  wire [30:0] n22838_o;
  wire [31:0] n22839_o;
  wire n22841_o;
  wire n22843_o;
  wire n22844_o;
  wire [5:0] n22846_o;
  wire [30:0] n22847_o;
  wire [31:0] n22848_o;
  wire n22850_o;
  wire n22852_o;
  wire n22853_o;
  wire [5:0] n22855_o;
  wire [30:0] n22856_o;
  wire [31:0] n22857_o;
  wire n22859_o;
  wire n22861_o;
  wire n22862_o;
  wire [5:0] n22864_o;
  wire [30:0] n22865_o;
  wire [31:0] n22866_o;
  wire n22868_o;
  wire n22870_o;
  wire n22871_o;
  wire [5:0] n22873_o;
  wire [30:0] n22874_o;
  wire [31:0] n22875_o;
  wire n22877_o;
  wire n22879_o;
  wire n22880_o;
  wire [5:0] n22882_o;
  wire [30:0] n22883_o;
  wire [31:0] n22884_o;
  wire n22886_o;
  wire n22888_o;
  wire n22889_o;
  wire [5:0] n22891_o;
  wire [30:0] n22892_o;
  wire [31:0] n22893_o;
  wire n22895_o;
  wire n22897_o;
  wire n22898_o;
  wire [5:0] n22900_o;
  wire [30:0] n22901_o;
  wire [31:0] n22902_o;
  wire n22904_o;
  wire n22906_o;
  wire n22907_o;
  wire [5:0] n22909_o;
  wire [30:0] n22910_o;
  wire [31:0] n22911_o;
  wire n22913_o;
  wire n22915_o;
  wire n22916_o;
  wire [5:0] n22918_o;
  wire [30:0] n22919_o;
  wire [31:0] n22920_o;
  wire n22922_o;
  wire n22924_o;
  wire n22925_o;
  wire [5:0] n22927_o;
  wire [30:0] n22928_o;
  wire [31:0] n22929_o;
  wire n22931_o;
  wire n22933_o;
  wire n22934_o;
  wire [5:0] n22936_o;
  wire [30:0] n22937_o;
  wire [31:0] n22938_o;
  wire n22940_o;
  wire n22942_o;
  wire n22943_o;
  wire [5:0] n22945_o;
  wire [30:0] n22946_o;
  wire [31:0] n22947_o;
  wire n22949_o;
  wire n22951_o;
  wire n22952_o;
  wire [5:0] n22954_o;
  wire [30:0] n22955_o;
  wire [31:0] n22956_o;
  wire n22958_o;
  wire n22960_o;
  wire n22961_o;
  wire [5:0] n22963_o;
  wire [30:0] n22964_o;
  wire [31:0] n22965_o;
  wire n22967_o;
  wire n22969_o;
  wire n22970_o;
  wire [5:0] n22972_o;
  wire [30:0] n22973_o;
  wire [31:0] n22974_o;
  wire n22976_o;
  wire n22978_o;
  wire n22979_o;
  wire [5:0] n22981_o;
  wire [30:0] n22982_o;
  wire [31:0] n22983_o;
  wire n22985_o;
  wire n22987_o;
  wire n22988_o;
  wire [5:0] n22990_o;
  wire [30:0] n22991_o;
  wire [31:0] n22992_o;
  wire n22994_o;
  wire n22996_o;
  wire n22997_o;
  wire [5:0] n22999_o;
  wire [30:0] n23000_o;
  wire [31:0] n23001_o;
  wire n23003_o;
  wire n23005_o;
  wire n23006_o;
  wire [5:0] n23008_o;
  wire [30:0] n23009_o;
  wire [31:0] n23010_o;
  wire n23012_o;
  wire n23014_o;
  wire n23015_o;
  wire [5:0] n23017_o;
  wire [30:0] n23018_o;
  wire [31:0] n23019_o;
  wire n23021_o;
  wire n23023_o;
  wire n23024_o;
  wire [5:0] n23026_o;
  wire [30:0] n23027_o;
  wire [31:0] n23028_o;
  wire n23030_o;
  wire n23032_o;
  wire n23033_o;
  wire n23034_o;
  wire [5:0] n23035_o;
  wire [30:0] n23036_o;
  wire [31:0] n23037_o;
  wire n23039_o;
  wire n23041_o;
  wire [43:0] n23042_o;
  wire [99:0] n23085_o;
  wire [66:0] n23086_o;
  wire [7:0] n23087_o;
  wire [7:0] n23088_o;
  wire [7:0] n23089_o;
  wire [7:0] n23090_o;
  wire [7:0] n23091_o;
  wire [7:0] n23092_o;
  wire [7:0] n23093_o;
  wire [7:0] n23094_o;
  wire [3:0] n23095_o;
  wire n23096_o;
  wire n23097_o;
  wire [63:0] n23098_o;
  wire n23099_o;
  wire [63:0] n23100_o;
  wire n23101_o;
  wire n23102_o;
  wire [63:0] n23103_o;
  wire [1:0] n23104_o;
  wire [2:0] n23106_o;
  wire [2:0] n23107_o;
  wire [5:0] n23108_o;
  wire [4:0] n23109_o;
  wire [5:0] n23111_o;
  wire [4:0] n23112_o;
  wire [47:0] n23113_o;
  wire [55:0] n23115_o;
  wire n23116_o;
  wire [63:0] n23117_o;
  wire n23118_o;
  wire n23119_o;
  wire n23120_o;
  wire n23121_o;
  wire n23122_o;
  wire n23123_o;
  wire n23124_o;
  wire n23125_o;
  wire n23126_o;
  wire n23127_o;
  wire n23128_o;
  wire n23129_o;
  wire n23130_o;
  wire n23131_o;
  wire n23132_o;
  wire n23133_o;
  wire n23134_o;
  wire n23135_o;
  wire n23136_o;
  wire n23140_o;
  wire n23141_o;
  wire n23142_o;
  wire n23143_o;
  wire n23144_o;
  wire n23145_o;
  wire n23148_o;
  wire n23149_o;
  wire n23151_o;
  wire [4:0] n23152_o;
  wire [5:0] n23154_o;
  wire n23157_o;
  wire [3:0] n23161_o;
  wire n23162_o;
  wire [3:0] n23163_o;
  wire [5:0] n23164_o;
  wire n23165_o;
  wire [3:0] n23166_o;
  wire [5:0] n23167_o;
  wire n23168_o;
  wire n23169_o;
  wire n23170_o;
  wire [3:0] n23171_o;
  wire n23173_o;
  wire n23175_o;
  wire n23177_o;
  wire [5:0] n23178_o;
  wire n23179_o;
  wire [68:0] n23180_o;
  wire [6:0] n23181_o;
  wire [68:0] n23182_o;
  wire [3:0] n23184_o;
  wire [3:0] n23185_o;
  wire n23187_o;
  wire n23189_o;
  wire n23190_o;
  wire [6:0] n23191_o;
  wire n23193_o;
  wire n23194_o;
  wire n23195_o;
  wire n23196_o;
  wire [31:0] n23197_o;
  wire [63:0] n23198_o;
  wire [63:0] n23201_o;
  wire [63:0] n23202_o;
  wire [31:0] n23203_o;
  wire [31:0] n23204_o;
  wire n23205_o;
  wire n23206_o;
  wire n23207_o;
  wire n23208_o;
  wire n23209_o;
  wire [100:0] n23213_o;
  wire n23214_o;
  wire n23215_o;
  wire n23216_o;
  wire [95:0] n23217_o;
  wire [100:0] n23218_o;
  wire [100:0] n23219_o;
  wire n23220_o;
  wire n23221_o;
  wire n23222_o;
  wire n23223_o;
  wire n23224_o;
  wire n23225_o;
  wire [67:0] n23226_o;
  wire [67:0] n23227_o;
  wire [67:0] n23228_o;
  wire [5:0] n23229_o;
  wire [5:0] n23230_o;
  wire [5:0] n23231_o;
  wire n23233_o;
  wire n23236_o;
  wire n23237_o;
  wire [3:0] n23239_o;
  wire [3:0] n23240_o;
  wire n23242_o;
  wire n23245_o;
  wire n23246_o;
  wire [63:0] n23247_o;
  wire [64:0] n23250_o;
  wire [3:0] n23251_o;
  wire [3:0] n23252_o;
  wire [64:0] n23253_o;
  wire [64:0] n23254_o;
  wire n23256_o;
  wire [4:0] n23257_o;
  wire [5:0] n23259_o;
  wire n23262_o;
  wire n23265_o;
  wire n23266_o;
  wire n23267_o;
  wire [63:0] n23268_o;
  wire [63:0] n23270_o;
  wire [64:0] n23272_o;
  wire [64:0] n23273_o;
  wire [64:0] n23274_o;
  wire [64:0] n23275_o;
  wire [64:0] n23276_o;
  wire [64:0] n23277_o;
  wire [63:0] n23278_o;
  wire [1:0] n23279_o;
  wire [2:0] n23281_o;
  wire [63:0] n23282_o;
  wire [2:0] n23283_o;
  wire [5:0] n23284_o;
  wire [63:0] n23285_o;
  wire [4:0] n23286_o;
  wire [5:0] n23288_o;
  wire [4:0] n23289_o;
  wire [63:0] n23290_o;
  wire [47:0] n23291_o;
  wire [55:0] n23293_o;
  wire n23295_o;
  wire [3:0] n23299_o;
  wire n23300_o;
  wire [196:0] n23301_o;
  wire [3:0] n23302_o;
  wire [3:0] n23303_o;
  wire [196:0] n23304_o;
  wire [196:0] n23305_o;
  wire n23306_o;
  wire n23309_o;
  wire [3:0] n23312_o;
  wire n23313_o;
  wire n23315_o;
  wire [4:0] n23316_o;
  wire [5:0] n23318_o;
  wire [5:0] n23319_o;
  wire [5:0] n23321_o;
  wire [5:0] n23322_o;
  wire [30:0] n23323_o;
  wire [30:0] n23324_o;
  wire [30:0] n23325_o;
  wire [30:0] n23326_o;
  wire n23327_o;
  wire n23328_o;
  wire n23329_o;
  wire n23330_o;
  wire n23331_o;
  wire n23335_o;
  wire n23337_o;
  wire n23338_o;
  wire [5:0] n23339_o;
  wire [5:0] n23341_o;
  wire n23342_o;
  wire n23343_o;
  wire [3:0] n23347_o;
  wire n23348_o;
  wire [3:0] n23349_o;
  wire n23350_o;
  wire n23351_o;
  wire n23353_o;
  wire n23356_o;
  wire n23357_o;
  wire [63:0] n23358_o;
  wire [63:0] n23359_o;
  wire n23360_o;
  wire [63:0] n23361_o;
  wire n23362_o;
  wire n23363_o;
  wire [63:0] n23364_o;
  wire n23365_o;
  wire n23366_o;
  wire n23367_o;
  wire n23368_o;
  wire n23369_o;
  wire [63:0] n23370_o;
  wire n23371_o;
  wire [63:0] n23372_o;
  wire n23373_o;
  wire n23374_o;
  wire n23375_o;
  wire n23376_o;
  wire n23377_o;
  wire [63:0] n23378_o;
  wire n23379_o;
  wire [63:0] n23380_o;
  wire n23381_o;
  wire n23382_o;
  wire n23383_o;
  wire n23384_o;
  wire n23386_o;
  wire [63:0] n23388_o;
  wire n23389_o;
  wire [63:0] n23390_o;
  wire n23391_o;
  wire n23392_o;
  wire n23393_o;
  wire n23394_o;
  wire n23395_o;
  wire n23396_o;
  wire n23399_o;
  wire [1:0] n23400_o;
  wire [3:0] n23401_o;
  wire [1:0] n23402_o;
  wire [1:0] n23403_o;
  wire [63:0] n23404_o;
  wire [4:0] n23405_o;
  wire [5:0] n23407_o;
  wire n23409_o;
  wire n23411_o;
  wire n23412_o;
  wire [5:0] n23413_o;
  wire n23414_o;
  wire n23415_o;
  wire [261:0] n23418_o;
  wire [501:0] n23419_o;
  wire [5:0] n23420_o;
  wire [5:0] n23421_o;
  wire [4:0] n23422_o;
  wire [63:0] n23423_o;
  wire [47:0] n23424_o;
  wire [55:0] n23426_o;
  wire [66:0] n23428_o;
  wire [3:0] n23429_o;
  wire [66:0] n23430_o;
  wire [66:0] n23431_o;
  wire n23432_o;
  wire [3:0] n23433_o;
  wire [66:0] n23434_o;
  wire [66:0] n23435_o;
  wire n23436_o;
  wire [1:0] n23437_o;
  wire [1:0] n23438_o;
  wire [3:0] n23444_o;
  wire [66:0] n23445_o;
  wire [66:0] n23446_o;
  wire n23447_o;
  wire n23448_o;
  wire [1:0] n23449_o;
  wire [1:0] n23450_o;
  wire [132:0] n23454_o;
  wire [3:0] n23455_o;
  wire [3:0] n23456_o;
  wire [130:0] n23457_o;
  wire [132:0] n23458_o;
  wire [1:0] n23460_o;
  wire [1:0] n23461_o;
  wire n23465_o;
  wire [3:0] n23468_o;
  wire n23469_o;
  wire n23470_o;
  wire n23471_o;
  wire n23472_o;
  wire [131:0] n23473_o;
  wire [131:0] n23474_o;
  wire [131:0] n23475_o;
  wire n23477_o;
  wire n23478_o;
  wire n23479_o;
  wire [3:0] n23482_o;
  wire n23485_o;
  wire n23488_o;
  wire n23490_o;
  wire n23493_o;
  wire [12:0] n23494_o;
  wire [67:0] n23495_o;
  reg [67:0] n23497_o;
  wire [96:0] n23498_o;
  wire [95:0] n23499_o;
  wire [96:0] n23500_o;
  reg [96:0] n23502_o;
  wire [3:0] n23503_o;
  reg [3:0] n23505_o;
  wire [63:0] n23506_o;
  wire [63:0] n23507_o;
  reg [63:0] n23509_o;
  wire n23510_o;
  wire n23511_o;
  reg n23513_o;
  wire [63:0] n23514_o;
  wire [63:0] n23515_o;
  reg [63:0] n23517_o;
  wire n23518_o;
  wire n23519_o;
  reg n23521_o;
  wire [63:0] n23522_o;
  wire [63:0] n23523_o;
  reg [63:0] n23525_o;
  wire n23526_o;
  wire n23527_o;
  reg n23529_o;
  wire [5:0] n23530_o;
  wire [5:0] n23531_o;
  wire [5:0] n23532_o;
  reg [5:0] n23534_o;
  wire [4:0] n23535_o;
  wire [4:0] n23536_o;
  wire [4:0] n23537_o;
  reg [4:0] n23539_o;
  wire [55:0] n23540_o;
  wire [55:0] n23541_o;
  wire [55:0] n23542_o;
  reg [55:0] n23544_o;
  wire [63:0] n23545_o;
  wire [63:0] n23546_o;
  reg [63:0] n23548_o;
  wire n23549_o;
  reg n23551_o;
  reg n23553_o;
  reg n23555_o;
  wire [1:0] n23556_o;
  reg [1:0] n23558_o;
  reg n23575_o;
  reg n23580_o;
  reg n23584_o;
  reg n23589_o;
  reg n23594_o;
  reg n23599_o;
  wire [501:0] n23615_o;
  wire [3:0] n23616_o;
  wire n23618_o;
  wire [501:0] n23619_o;
  wire [3:0] n23620_o;
  wire n23622_o;
  wire n23623_o;
  wire n23624_o;
  wire n23625_o;
  wire [501:0] n23626_o;
  wire n23627_o;
  wire [501:0] n23628_o;
  wire n23629_o;
  wire n23630_o;
  wire [501:0] n23631_o;
  wire n23632_o;
  wire n23633_o;
  wire [501:0] n23634_o;
  wire n23635_o;
  wire n23636_o;
  wire [501:0] n23637_o;
  wire n23638_o;
  wire n23639_o;
  wire [501:0] n23640_o;
  wire n23641_o;
  wire n23642_o;
  wire [1:0] n23643_o;
  wire [1:0] n23644_o;
  wire [1:0] n23645_o;
  wire n23646_o;
  wire [31:0] n23647_o;
  wire [31:0] n23649_o;
  wire [19:0] n23650_o;
  wire [27:0] n23652_o;
  wire [23:0] n23653_o;
  wire [23:0] n23654_o;
  wire [23:0] n23655_o;
  wire [23:0] n23656_o;
  wire [23:0] n23657_o;
  wire [23:0] n23658_o;
  wire [23:0] n23659_o;
  wire [23:0] n23660_o;
  wire [51:0] n23661_o;
  wire [7:0] n23662_o;
  wire [59:0] n23663_o;
  wire [63:0] n23665_o;
  wire [36:0] n23666_o;
  wire [44:0] n23668_o;
  wire [15:0] n23669_o;
  wire [15:0] n23670_o;
  wire [15:0] n23671_o;
  wire [15:0] n23672_o;
  wire [15:0] n23673_o;
  wire [60:0] n23674_o;
  wire [63:0] n23676_o;
  wire [43:0] n23677_o;
  wire [43:0] n23678_o;
  wire [43:0] n23679_o;
  wire [43:0] n23680_o;
  wire [43:0] n23681_o;
  wire [43:0] n23682_o;
  wire [51:0] n23684_o;
  wire [11:0] n23685_o;
  wire [63:0] n23686_o;
  wire [501:0] n23687_o;
  wire [63:0] n23688_o;
  wire [51:0] n23689_o;
  wire [63:0] n23691_o;
  wire [43:0] n23692_o;
  wire [51:0] n23694_o;
  wire [63:0] n23696_o;
  wire [63:0] n23697_o;
  wire [63:0] n23698_o;
  wire [63:0] n23700_o;
  wire [63:0] n23701_o;
  wire [63:0] n23703_o;
  wire [63:0] n23704_o;
  wire n23705_o;
  wire n23706_o;
  wire n23707_o;
  wire n23708_o;
  wire n23709_o;
  wire n23710_o;
  wire n23711_o;
  wire n23712_o;
  wire n23713_o;
  reg [501:0] n23721_q;
  wire [70:0] n23722_o;
  wire [131:0] n23723_o;
  wire [130:0] n23724_o;
  assign l_out_done = n22423_o;
  assign l_out_err = n22424_o;
  assign l_out_invalid = n22425_o;
  assign l_out_badtree = n22426_o;
  assign l_out_segerr = n22427_o;
  assign l_out_perm_error = n22428_o;
  assign l_out_rc_error = n22429_o;
  assign l_out_sprval = n22430_o;
  assign d_out_valid = n22432_o;
  assign d_out_tlbie = n22433_o;
  assign d_out_doall = n22434_o;
  assign d_out_tlbld = n22435_o;
  assign d_out_addr = n22436_o;
  assign d_out_pte = n22437_o;
  assign i_out_tlbld = n22440_o;
  assign i_out_tlbie = n22441_o;
  assign i_out_doall = n22442_o;
  assign i_out_addr = n22443_o;
  assign i_out_pte = n22444_o;
  /* loadstore1.vhdl:685:63  */
  assign n22421_o = {l_in_rs, l_in_addr, l_in_sprn, l_in_priv, l_in_load, l_in_iside, l_in_mtspr, l_in_slbia, l_in_tlbie, l_in_valid};
  assign n22423_o = n23722_o[0];
  assign n22424_o = n23722_o[1];
  assign n22425_o = n23722_o[2];
  assign n22426_o = n23722_o[3];
  /* loadstore1.vhdl:645:5  */
  assign n22427_o = n23722_o[4];
  /* loadstore1.vhdl:663:18  */
  assign n22428_o = n23722_o[5];
  assign n22429_o = n23722_o[6];
  /* loadstore1.vhdl:662:18  */
  assign n22430_o = n23722_o[70:7];
  /* loadstore1.vhdl:661:18  */
  assign n22432_o = n23723_o[0];
  assign n22433_o = n23723_o[1];
  /* loadstore1.vhdl:660:18  */
  assign n22434_o = n23723_o[2];
  assign n22435_o = n23723_o[3];
  /* loadstore1.vhdl:659:18  */
  assign n22436_o = n23723_o[67:4];
  assign n22437_o = n23723_o[131:68];
  /* loadstore1.vhdl:658:18  */
  assign n22438_o = {d_in_data, d_in_err, d_in_done, d_in_stall};
  /* loadstore1.vhdl:657:18  */
  assign n22440_o = n23724_o[0];
  assign n22441_o = n23724_o[1];
  /* loadstore1.vhdl:656:18  */
  assign n22442_o = n23724_o[2];
  assign n22443_o = n23724_o[66:3];
  /* loadstore1.vhdl:655:18  */
  assign n22444_o = n23724_o[130:67];
  /* mmu.vhdl:76:12  */
  assign r = n23721_q; // (signal)
  /* mmu.vhdl:76:15  */
  assign rin = n23687_o; // (signal)
  /* mmu.vhdl:78:12  */
  assign addrsh = n22539_o; // (signal)
  /* mmu.vhdl:79:12  */
  assign mask = n22642_o; // (signal)
  /* mmu.vhdl:80:12  */
  assign finalmask = n23042_o; // (signal)
  /* mmu.vhdl:85:23  */
  assign n22445_o = r[132:69];
  /* mmu.vhdl:85:42  */
  assign n22446_o = n22421_o[15];
  /* mmu.vhdl:85:28  */
  assign n22447_o = n22446_o ? n22445_o : n22450_o;
  /* mmu.vhdl:85:73  */
  assign n22448_o = r[164:133];
  /* mmu.vhdl:85:69  */
  assign n22450_o = {32'b00000000000000000000000000000000, n22448_o};
  /* loadstore1.vhdl:594:32  */
  assign n22469_o = {4'b0000, 32'b00000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000};
  assign n22470_o = rin[0];
  /* mmu.vhdl:90:13  */
  assign n22471_o = rst ? 1'b0 : n22470_o;
  /* loadstore1.vhdl:594:18  */
  assign n22472_o = rin[68:1];
  /* loadstore1.vhdl:595:71  */
  assign n22473_o = r[68:1];
  /* mmu.vhdl:90:13  */
  assign n22474_o = rst ? n22473_o : n22472_o;
  /* loadstore1.vhdl:594:32  */
  assign n22475_o = rin[168:69];
  /* mmu.vhdl:90:13  */
  assign n22476_o = rst ? n22469_o : n22475_o;
  /* loadstore1.vhdl:594:32  */
  assign n22477_o = rin[234:169];
  /* loadstore1.vhdl:594:18  */
  assign n22478_o = r[234:169];
  /* mmu.vhdl:90:13  */
  assign n22479_o = rst ? n22478_o : n22477_o;
  assign n22480_o = rin[235];
  /* mmu.vhdl:90:13  */
  assign n22481_o = rst ? 1'b0 : n22480_o;
  assign n22482_o = rin[299:236];
  /* loadstore1.vhdl:594:32  */
  assign n22483_o = r[299:236];
  /* mmu.vhdl:90:13  */
  assign n22484_o = rst ? n22483_o : n22482_o;
  /* loadstore1.vhdl:595:71  */
  assign n22485_o = rin[300];
  /* mmu.vhdl:90:13  */
  assign n22486_o = rst ? 1'b0 : n22485_o;
  /* loadstore1.vhdl:594:32  */
  assign n22487_o = rin[364:301];
  assign n22488_o = r[364:301];
  /* mmu.vhdl:90:13  */
  assign n22489_o = rst ? n22488_o : n22487_o;
  /* loadstore1.vhdl:594:18  */
  assign n22490_o = rin[365];
  /* mmu.vhdl:90:13  */
  assign n22491_o = rst ? 1'b0 : n22490_o;
  assign n22492_o = rin[501:366];
  /* loadstore1.vhdl:594:32  */
  assign n22493_o = r[501:366];
  /* mmu.vhdl:90:13  */
  assign n22494_o = rst ? n22493_o : n22492_o;
  /* loadstore1.vhdl:594:32  */
  assign n22495_o = {n22494_o, n22491_o, n22489_o, n22486_o, n22484_o, n22481_o, n22479_o, n22476_o, n22474_o, n22471_o};
  /* mmu.vhdl:129:21  */
  assign n22502_o = r[371:370];
  /* mmu.vhdl:131:30  */
  assign n22503_o = r[46:16];
  /* mmu.vhdl:130:13  */
  assign n22505_o = n22502_o == 2'b00;
  /* mmu.vhdl:133:30  */
  assign n22506_o = r[62:32];
  /* mmu.vhdl:132:13  */
  assign n22508_o = n22502_o == 2'b01;
  /* mmu.vhdl:135:48  */
  assign n22509_o = r[65:48];
  /* mmu.vhdl:135:40  */
  assign n22511_o = {13'b0000000000000, n22509_o};
  /* loadstore1.vhdl:579:5  */
  assign n22512_o = {n22508_o, n22505_o};
  /* mmu.vhdl:129:9  */
  always @*
    case (n22512_o)
      2'b10: n22513_o = n22506_o;
      2'b01: n22513_o = n22503_o;
      default: n22513_o = n22511_o;
    endcase
  /* mmu.vhdl:137:21  */
  assign n22514_o = r[369:368];
  /* mmu.vhdl:139:27  */
  assign n22515_o = n22513_o[18:0];
  /* mmu.vhdl:138:13  */
  assign n22517_o = n22514_o == 2'b00;
  /* mmu.vhdl:141:27  */
  assign n22518_o = n22513_o[22:4];
  /* mmu.vhdl:140:13  */
  assign n22520_o = n22514_o == 2'b01;
  /* mmu.vhdl:143:27  */
  assign n22521_o = n22513_o[26:8];
  /* mmu.vhdl:142:13  */
  assign n22523_o = n22514_o == 2'b10;
  /* mmu.vhdl:145:27  */
  assign n22524_o = n22513_o[30:12];
  assign n22525_o = {n22523_o, n22520_o, n22517_o};
  /* mmu.vhdl:137:9  */
  always @*
    case (n22525_o)
      3'b100: n22526_o = n22521_o;
      3'b010: n22526_o = n22518_o;
      3'b001: n22526_o = n22515_o;
      default: n22526_o = n22524_o;
    endcase
  /* mmu.vhdl:147:21  */
  assign n22527_o = r[367:366];
  /* mmu.vhdl:149:30  */
  assign n22528_o = n22526_o[15:0];
  /* mmu.vhdl:148:13  */
  assign n22530_o = n22527_o == 2'b00;
  /* mmu.vhdl:151:30  */
  assign n22531_o = n22526_o[16:1];
  /* mmu.vhdl:150:13  */
  assign n22533_o = n22527_o == 2'b01;
  /* mmu.vhdl:153:30  */
  assign n22534_o = n22526_o[17:2];
  /* mmu.vhdl:152:13  */
  assign n22536_o = n22527_o == 2'b10;
  /* mmu.vhdl:155:30  */
  assign n22537_o = n22526_o[18:3];
  assign n22538_o = {n22536_o, n22533_o, n22530_o};
  /* mmu.vhdl:147:9  */
  always @*
    case (n22538_o)
      3'b100: n22539_o = n22534_o;
      3'b010: n22539_o = n22531_o;
      3'b001: n22539_o = n22528_o;
      default: n22539_o = n22537_o;
    endcase
  /* mmu.vhdl:167:33  */
  assign n22543_o = r[376:372];
  /* mmu.vhdl:167:20  */
  assign n22544_o = {26'b0, n22543_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22545_o = {1'b0, n22544_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22547_o = $signed(32'b00000000000000000000000000000101) < $signed(n22545_o);
  /* mmu.vhdl:167:13  */
  assign n22550_o = n22547_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:631:18  */
  assign n22553_o = n22551_o[4:0];
  /* mmu.vhdl:167:33  */
  assign n22554_o = r[376:372];
  /* mmu.vhdl:167:20  */
  assign n22555_o = {26'b0, n22554_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22556_o = {1'b0, n22555_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22558_o = $signed(32'b00000000000000000000000000000110) < $signed(n22556_o);
  /* fpu.vhdl:635:18  */
  assign n22560_o = n22551_o[6];
  /* mmu.vhdl:167:13  */
  assign n22561_o = n22558_o ? 1'b1 : n22560_o;
  /* mmu.vhdl:167:33  */
  assign n22563_o = r[376:372];
  /* mmu.vhdl:167:20  */
  assign n22564_o = {26'b0, n22563_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22565_o = {1'b0, n22564_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22567_o = $signed(32'b00000000000000000000000000000111) < $signed(n22565_o);
  /* loadstore1.vhdl:199:18  */
  assign n22569_o = n22551_o[7];
  /* mmu.vhdl:167:13  */
  assign n22570_o = n22567_o ? 1'b1 : n22569_o;
  /* mmu.vhdl:167:33  */
  assign n22572_o = r[376:372];
  /* mmu.vhdl:167:20  */
  assign n22573_o = {26'b0, n22572_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22574_o = {1'b0, n22573_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22576_o = $signed(32'b00000000000000000000000000001000) < $signed(n22574_o);
  /* fpu.vhdl:997:17  */
  assign n22578_o = n22551_o[8];
  /* mmu.vhdl:167:13  */
  assign n22579_o = n22576_o ? 1'b1 : n22578_o;
  /* mmu.vhdl:167:33  */
  assign n22581_o = r[376:372];
  /* mmu.vhdl:167:20  */
  assign n22582_o = {26'b0, n22581_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22583_o = {1'b0, n22582_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22585_o = $signed(32'b00000000000000000000000000001001) < $signed(n22583_o);
  assign n22587_o = n22551_o[9];
  /* mmu.vhdl:167:13  */
  assign n22588_o = n22585_o ? 1'b1 : n22587_o;
  /* mmu.vhdl:167:33  */
  assign n22590_o = r[376:372];
  /* mmu.vhdl:167:20  */
  assign n22591_o = {26'b0, n22590_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22592_o = {1'b0, n22591_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22594_o = $signed(32'b00000000000000000000000000001010) < $signed(n22592_o);
  /* loadstore1.vhdl:377:47  */
  assign n22596_o = n22551_o[10];
  /* mmu.vhdl:167:13  */
  assign n22597_o = n22594_o ? 1'b1 : n22596_o;
  /* mmu.vhdl:167:33  */
  assign n22599_o = r[376:372];
  /* mmu.vhdl:167:20  */
  assign n22600_o = {26'b0, n22599_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22601_o = {1'b0, n22600_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22603_o = $signed(32'b00000000000000000000000000001011) < $signed(n22601_o);
  /* loadstore1.vhdl:373:18  */
  assign n22605_o = n22551_o[11];
  /* mmu.vhdl:167:13  */
  assign n22606_o = n22603_o ? 1'b1 : n22605_o;
  /* mmu.vhdl:167:33  */
  assign n22608_o = r[376:372];
  /* mmu.vhdl:167:20  */
  assign n22609_o = {26'b0, n22608_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22610_o = {1'b0, n22609_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22612_o = $signed(32'b00000000000000000000000000001100) < $signed(n22610_o);
  assign n22614_o = n22551_o[12];
  /* mmu.vhdl:167:13  */
  assign n22615_o = n22612_o ? 1'b1 : n22614_o;
  /* mmu.vhdl:167:33  */
  assign n22617_o = r[376:372];
  /* mmu.vhdl:167:20  */
  assign n22618_o = {26'b0, n22617_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22619_o = {1'b0, n22618_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22621_o = $signed(32'b00000000000000000000000000001101) < $signed(n22619_o);
  assign n22623_o = n22551_o[13];
  /* mmu.vhdl:167:13  */
  assign n22624_o = n22621_o ? 1'b1 : n22623_o;
  /* mmu.vhdl:167:33  */
  assign n22626_o = r[376:372];
  /* mmu.vhdl:167:20  */
  assign n22627_o = {26'b0, n22626_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22628_o = {1'b0, n22627_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22630_o = $signed(32'b00000000000000000000000000001110) < $signed(n22628_o);
  /* loadstore1.vhdl:338:22  */
  assign n22632_o = n22551_o[14];
  /* mmu.vhdl:167:13  */
  assign n22633_o = n22630_o ? 1'b1 : n22632_o;
  /* loadstore1.vhdl:337:22  */
  assign n22634_o = n22551_o[15];
  /* mmu.vhdl:167:33  */
  assign n22635_o = r[376:372];
  /* mmu.vhdl:167:20  */
  assign n22636_o = {26'b0, n22635_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22637_o = {1'b0, n22636_o};  //  uext
  /* mmu.vhdl:167:18  */
  assign n22639_o = $signed(32'b00000000000000000000000000001111) < $signed(n22637_o);
  /* mmu.vhdl:167:13  */
  assign n22641_o = n22639_o ? 1'b1 : n22634_o;
  /* loadstore1.vhdl:333:22  */
  assign n22642_o = {n22641_o, n22633_o, n22624_o, n22615_o, n22606_o, n22597_o, n22588_o, n22579_o, n22570_o, n22561_o, n22550_o, n22553_o};
  /* mmu.vhdl:181:33  */
  assign n22647_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22648_o = {25'b0, n22647_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22649_o = {1'b0, n22648_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22651_o = $signed(32'b00000000000000000000000000000000) < $signed(n22649_o);
  /* mmu.vhdl:181:13  */
  assign n22654_o = n22651_o ? 1'b1 : 1'b0;
  /* mmu.vhdl:181:33  */
  assign n22657_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22658_o = {25'b0, n22657_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22659_o = {1'b0, n22658_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22661_o = $signed(32'b00000000000000000000000000000001) < $signed(n22659_o);
  assign n22663_o = n22655_o[1];
  /* mmu.vhdl:181:13  */
  assign n22664_o = n22661_o ? 1'b1 : n22663_o;
  /* mmu.vhdl:181:33  */
  assign n22666_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22667_o = {25'b0, n22666_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22668_o = {1'b0, n22667_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22670_o = $signed(32'b00000000000000000000000000000010) < $signed(n22668_o);
  /* loadstore1.vhdl:301:21  */
  assign n22672_o = n22655_o[2];
  /* mmu.vhdl:181:13  */
  assign n22673_o = n22670_o ? 1'b1 : n22672_o;
  /* mmu.vhdl:181:33  */
  assign n22675_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22676_o = {25'b0, n22675_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22677_o = {1'b0, n22676_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22679_o = $signed(32'b00000000000000000000000000000011) < $signed(n22677_o);
  assign n22681_o = n22655_o[3];
  /* mmu.vhdl:181:13  */
  assign n22682_o = n22679_o ? 1'b1 : n22681_o;
  /* mmu.vhdl:181:33  */
  assign n22684_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22685_o = {25'b0, n22684_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22686_o = {1'b0, n22685_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22688_o = $signed(32'b00000000000000000000000000000100) < $signed(n22686_o);
  assign n22690_o = n22655_o[4];
  /* mmu.vhdl:181:13  */
  assign n22691_o = n22688_o ? 1'b1 : n22690_o;
  /* mmu.vhdl:181:33  */
  assign n22693_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22694_o = {25'b0, n22693_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22695_o = {1'b0, n22694_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22697_o = $signed(32'b00000000000000000000000000000101) < $signed(n22695_o);
  assign n22699_o = n22655_o[5];
  /* mmu.vhdl:181:13  */
  assign n22700_o = n22697_o ? 1'b1 : n22699_o;
  /* mmu.vhdl:181:33  */
  assign n22702_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22703_o = {25'b0, n22702_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22704_o = {1'b0, n22703_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22706_o = $signed(32'b00000000000000000000000000000110) < $signed(n22704_o);
  assign n22708_o = n22655_o[6];
  /* mmu.vhdl:181:13  */
  assign n22709_o = n22706_o ? 1'b1 : n22708_o;
  /* mmu.vhdl:181:33  */
  assign n22711_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22712_o = {25'b0, n22711_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22713_o = {1'b0, n22712_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22715_o = $signed(32'b00000000000000000000000000000111) < $signed(n22713_o);
  assign n22717_o = n22655_o[7];
  /* mmu.vhdl:181:13  */
  assign n22718_o = n22715_o ? 1'b1 : n22717_o;
  /* mmu.vhdl:181:33  */
  assign n22720_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22721_o = {25'b0, n22720_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22722_o = {1'b0, n22721_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22724_o = $signed(32'b00000000000000000000000000001000) < $signed(n22722_o);
  assign n22726_o = n22655_o[8];
  /* mmu.vhdl:181:13  */
  assign n22727_o = n22724_o ? 1'b1 : n22726_o;
  /* mmu.vhdl:181:33  */
  assign n22729_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22730_o = {25'b0, n22729_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22731_o = {1'b0, n22730_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22733_o = $signed(32'b00000000000000000000000000001001) < $signed(n22731_o);
  assign n22735_o = n22655_o[9];
  /* mmu.vhdl:181:13  */
  assign n22736_o = n22733_o ? 1'b1 : n22735_o;
  /* mmu.vhdl:181:33  */
  assign n22738_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22739_o = {25'b0, n22738_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22740_o = {1'b0, n22739_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22742_o = $signed(32'b00000000000000000000000000001010) < $signed(n22740_o);
  assign n22744_o = n22655_o[10];
  /* mmu.vhdl:181:13  */
  assign n22745_o = n22742_o ? 1'b1 : n22744_o;
  /* mmu.vhdl:181:33  */
  assign n22747_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22748_o = {25'b0, n22747_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22749_o = {1'b0, n22748_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22751_o = $signed(32'b00000000000000000000000000001011) < $signed(n22749_o);
  assign n22753_o = n22655_o[11];
  /* mmu.vhdl:181:13  */
  assign n22754_o = n22751_o ? 1'b1 : n22753_o;
  /* mmu.vhdl:181:33  */
  assign n22756_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22757_o = {25'b0, n22756_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22758_o = {1'b0, n22757_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22760_o = $signed(32'b00000000000000000000000000001100) < $signed(n22758_o);
  assign n22762_o = n22655_o[12];
  /* mmu.vhdl:181:13  */
  assign n22763_o = n22760_o ? 1'b1 : n22762_o;
  /* mmu.vhdl:181:33  */
  assign n22765_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22766_o = {25'b0, n22765_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22767_o = {1'b0, n22766_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22769_o = $signed(32'b00000000000000000000000000001101) < $signed(n22767_o);
  assign n22771_o = n22655_o[13];
  /* mmu.vhdl:181:13  */
  assign n22772_o = n22769_o ? 1'b1 : n22771_o;
  /* mmu.vhdl:181:33  */
  assign n22774_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22775_o = {25'b0, n22774_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22776_o = {1'b0, n22775_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22778_o = $signed(32'b00000000000000000000000000001110) < $signed(n22776_o);
  assign n22780_o = n22655_o[14];
  /* mmu.vhdl:181:13  */
  assign n22781_o = n22778_o ? 1'b1 : n22780_o;
  /* mmu.vhdl:181:33  */
  assign n22783_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22784_o = {25'b0, n22783_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22785_o = {1'b0, n22784_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22787_o = $signed(32'b00000000000000000000000000001111) < $signed(n22785_o);
  assign n22789_o = n22655_o[15];
  /* mmu.vhdl:181:13  */
  assign n22790_o = n22787_o ? 1'b1 : n22789_o;
  /* mmu.vhdl:181:33  */
  assign n22792_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22793_o = {25'b0, n22792_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22794_o = {1'b0, n22793_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22796_o = $signed(32'b00000000000000000000000000010000) < $signed(n22794_o);
  assign n22798_o = n22655_o[16];
  /* mmu.vhdl:181:13  */
  assign n22799_o = n22796_o ? 1'b1 : n22798_o;
  /* mmu.vhdl:181:33  */
  assign n22801_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22802_o = {25'b0, n22801_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22803_o = {1'b0, n22802_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22805_o = $signed(32'b00000000000000000000000000010001) < $signed(n22803_o);
  assign n22807_o = n22655_o[17];
  /* mmu.vhdl:181:13  */
  assign n22808_o = n22805_o ? 1'b1 : n22807_o;
  /* mmu.vhdl:181:33  */
  assign n22810_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22811_o = {25'b0, n22810_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22812_o = {1'b0, n22811_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22814_o = $signed(32'b00000000000000000000000000010010) < $signed(n22812_o);
  assign n22816_o = n22655_o[18];
  /* mmu.vhdl:181:13  */
  assign n22817_o = n22814_o ? 1'b1 : n22816_o;
  /* mmu.vhdl:181:33  */
  assign n22819_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22820_o = {25'b0, n22819_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22821_o = {1'b0, n22820_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22823_o = $signed(32'b00000000000000000000000000010011) < $signed(n22821_o);
  assign n22825_o = n22655_o[19];
  /* mmu.vhdl:181:13  */
  assign n22826_o = n22823_o ? 1'b1 : n22825_o;
  /* mmu.vhdl:181:33  */
  assign n22828_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22829_o = {25'b0, n22828_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22830_o = {1'b0, n22829_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22832_o = $signed(32'b00000000000000000000000000010100) < $signed(n22830_o);
  assign n22834_o = n22655_o[20];
  /* mmu.vhdl:181:13  */
  assign n22835_o = n22832_o ? 1'b1 : n22834_o;
  /* mmu.vhdl:181:33  */
  assign n22837_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22838_o = {25'b0, n22837_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22839_o = {1'b0, n22838_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22841_o = $signed(32'b00000000000000000000000000010101) < $signed(n22839_o);
  assign n22843_o = n22655_o[21];
  /* mmu.vhdl:181:13  */
  assign n22844_o = n22841_o ? 1'b1 : n22843_o;
  /* mmu.vhdl:181:33  */
  assign n22846_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22847_o = {25'b0, n22846_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22848_o = {1'b0, n22847_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22850_o = $signed(32'b00000000000000000000000000010110) < $signed(n22848_o);
  assign n22852_o = n22655_o[22];
  /* mmu.vhdl:181:13  */
  assign n22853_o = n22850_o ? 1'b1 : n22852_o;
  /* mmu.vhdl:181:33  */
  assign n22855_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22856_o = {25'b0, n22855_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22857_o = {1'b0, n22856_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22859_o = $signed(32'b00000000000000000000000000010111) < $signed(n22857_o);
  assign n22861_o = n22655_o[23];
  /* mmu.vhdl:181:13  */
  assign n22862_o = n22859_o ? 1'b1 : n22861_o;
  /* mmu.vhdl:181:33  */
  assign n22864_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22865_o = {25'b0, n22864_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22866_o = {1'b0, n22865_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22868_o = $signed(32'b00000000000000000000000000011000) < $signed(n22866_o);
  assign n22870_o = n22655_o[24];
  /* mmu.vhdl:181:13  */
  assign n22871_o = n22868_o ? 1'b1 : n22870_o;
  /* mmu.vhdl:181:33  */
  assign n22873_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22874_o = {25'b0, n22873_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22875_o = {1'b0, n22874_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22877_o = $signed(32'b00000000000000000000000000011001) < $signed(n22875_o);
  assign n22879_o = n22655_o[25];
  /* mmu.vhdl:181:13  */
  assign n22880_o = n22877_o ? 1'b1 : n22879_o;
  /* mmu.vhdl:181:33  */
  assign n22882_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22883_o = {25'b0, n22882_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22884_o = {1'b0, n22883_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22886_o = $signed(32'b00000000000000000000000000011010) < $signed(n22884_o);
  assign n22888_o = n22655_o[26];
  /* mmu.vhdl:181:13  */
  assign n22889_o = n22886_o ? 1'b1 : n22888_o;
  /* mmu.vhdl:181:33  */
  assign n22891_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22892_o = {25'b0, n22891_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22893_o = {1'b0, n22892_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22895_o = $signed(32'b00000000000000000000000000011011) < $signed(n22893_o);
  assign n22897_o = n22655_o[27];
  /* mmu.vhdl:181:13  */
  assign n22898_o = n22895_o ? 1'b1 : n22897_o;
  /* mmu.vhdl:181:33  */
  assign n22900_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22901_o = {25'b0, n22900_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22902_o = {1'b0, n22901_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22904_o = $signed(32'b00000000000000000000000000011100) < $signed(n22902_o);
  assign n22906_o = n22655_o[28];
  /* mmu.vhdl:181:13  */
  assign n22907_o = n22904_o ? 1'b1 : n22906_o;
  /* mmu.vhdl:181:33  */
  assign n22909_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22910_o = {25'b0, n22909_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22911_o = {1'b0, n22910_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22913_o = $signed(32'b00000000000000000000000000011101) < $signed(n22911_o);
  assign n22915_o = n22655_o[29];
  /* mmu.vhdl:181:13  */
  assign n22916_o = n22913_o ? 1'b1 : n22915_o;
  /* mmu.vhdl:181:33  */
  assign n22918_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22919_o = {25'b0, n22918_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22920_o = {1'b0, n22919_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22922_o = $signed(32'b00000000000000000000000000011110) < $signed(n22920_o);
  assign n22924_o = n22655_o[30];
  /* mmu.vhdl:181:13  */
  assign n22925_o = n22922_o ? 1'b1 : n22924_o;
  /* mmu.vhdl:181:33  */
  assign n22927_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22928_o = {25'b0, n22927_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22929_o = {1'b0, n22928_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22931_o = $signed(32'b00000000000000000000000000011111) < $signed(n22929_o);
  assign n22933_o = n22655_o[31];
  /* mmu.vhdl:181:13  */
  assign n22934_o = n22931_o ? 1'b1 : n22933_o;
  /* mmu.vhdl:181:33  */
  assign n22936_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22937_o = {25'b0, n22936_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22938_o = {1'b0, n22937_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22940_o = $signed(32'b00000000000000000000000000100000) < $signed(n22938_o);
  assign n22942_o = n22655_o[32];
  /* mmu.vhdl:181:13  */
  assign n22943_o = n22940_o ? 1'b1 : n22942_o;
  /* mmu.vhdl:181:33  */
  assign n22945_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22946_o = {25'b0, n22945_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22947_o = {1'b0, n22946_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22949_o = $signed(32'b00000000000000000000000000100001) < $signed(n22947_o);
  assign n22951_o = n22655_o[33];
  /* mmu.vhdl:181:13  */
  assign n22952_o = n22949_o ? 1'b1 : n22951_o;
  /* mmu.vhdl:181:33  */
  assign n22954_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22955_o = {25'b0, n22954_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22956_o = {1'b0, n22955_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22958_o = $signed(32'b00000000000000000000000000100010) < $signed(n22956_o);
  assign n22960_o = n22655_o[34];
  /* mmu.vhdl:181:13  */
  assign n22961_o = n22958_o ? 1'b1 : n22960_o;
  /* mmu.vhdl:181:33  */
  assign n22963_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22964_o = {25'b0, n22963_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22965_o = {1'b0, n22964_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22967_o = $signed(32'b00000000000000000000000000100011) < $signed(n22965_o);
  assign n22969_o = n22655_o[35];
  /* mmu.vhdl:181:13  */
  assign n22970_o = n22967_o ? 1'b1 : n22969_o;
  /* mmu.vhdl:181:33  */
  assign n22972_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22973_o = {25'b0, n22972_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22974_o = {1'b0, n22973_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22976_o = $signed(32'b00000000000000000000000000100100) < $signed(n22974_o);
  assign n22978_o = n22655_o[36];
  /* mmu.vhdl:181:13  */
  assign n22979_o = n22976_o ? 1'b1 : n22978_o;
  /* mmu.vhdl:181:33  */
  assign n22981_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22982_o = {25'b0, n22981_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22983_o = {1'b0, n22982_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22985_o = $signed(32'b00000000000000000000000000100101) < $signed(n22983_o);
  assign n22987_o = n22655_o[37];
  /* mmu.vhdl:181:13  */
  assign n22988_o = n22985_o ? 1'b1 : n22987_o;
  /* mmu.vhdl:181:33  */
  assign n22990_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n22991_o = {25'b0, n22990_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22992_o = {1'b0, n22991_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n22994_o = $signed(32'b00000000000000000000000000100110) < $signed(n22992_o);
  assign n22996_o = n22655_o[38];
  /* mmu.vhdl:181:13  */
  assign n22997_o = n22994_o ? 1'b1 : n22996_o;
  /* mmu.vhdl:181:33  */
  assign n22999_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n23000_o = {25'b0, n22999_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n23001_o = {1'b0, n23000_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n23003_o = $signed(32'b00000000000000000000000000100111) < $signed(n23001_o);
  assign n23005_o = n22655_o[39];
  /* mmu.vhdl:181:13  */
  assign n23006_o = n23003_o ? 1'b1 : n23005_o;
  /* mmu.vhdl:181:33  */
  assign n23008_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n23009_o = {25'b0, n23008_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n23010_o = {1'b0, n23009_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n23012_o = $signed(32'b00000000000000000000000000101000) < $signed(n23010_o);
  assign n23014_o = n22655_o[40];
  /* mmu.vhdl:181:13  */
  assign n23015_o = n23012_o ? 1'b1 : n23014_o;
  /* mmu.vhdl:181:33  */
  assign n23017_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n23018_o = {25'b0, n23017_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n23019_o = {1'b0, n23018_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n23021_o = $signed(32'b00000000000000000000000000101001) < $signed(n23019_o);
  assign n23023_o = n22655_o[41];
  /* mmu.vhdl:181:13  */
  assign n23024_o = n23021_o ? 1'b1 : n23023_o;
  /* mmu.vhdl:181:33  */
  assign n23026_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n23027_o = {25'b0, n23026_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n23028_o = {1'b0, n23027_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n23030_o = $signed(32'b00000000000000000000000000101010) < $signed(n23028_o);
  assign n23032_o = n22655_o[42];
  /* mmu.vhdl:181:13  */
  assign n23033_o = n23030_o ? 1'b1 : n23032_o;
  assign n23034_o = n22655_o[43];
  /* mmu.vhdl:181:33  */
  assign n23035_o = r[371:366];
  /* mmu.vhdl:181:20  */
  assign n23036_o = {25'b0, n23035_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n23037_o = {1'b0, n23036_o};  //  uext
  /* mmu.vhdl:181:18  */
  assign n23039_o = $signed(32'b00000000000000000000000000101011) < $signed(n23037_o);
  /* mmu.vhdl:181:13  */
  assign n23041_o = n23039_o ? 1'b1 : n23034_o;
  assign n23042_o = {n23041_o, n23033_o, n23024_o, n23015_o, n23006_o, n22997_o, n22988_o, n22979_o, n22970_o, n22961_o, n22952_o, n22943_o, n22934_o, n22925_o, n22916_o, n22907_o, n22898_o, n22889_o, n22880_o, n22871_o, n22862_o, n22853_o, n22844_o, n22835_o, n22826_o, n22817_o, n22808_o, n22799_o, n22790_o, n22781_o, n22772_o, n22763_o, n22754_o, n22745_o, n22736_o, n22727_o, n22718_o, n22709_o, n22700_o, n22691_o, n22682_o, n22673_o, n22664_o, n22654_o};
  assign n23085_o = r[168:69];
  assign n23086_o = r[67:1];
  /* mmu.vhdl:231:54  */
  assign n23087_o = n22438_o[66:59];
  /* mmu.vhdl:231:54  */
  assign n23088_o = n22438_o[58:51];
  /* mmu.vhdl:231:54  */
  assign n23089_o = n22438_o[50:43];
  /* mmu.vhdl:231:54  */
  assign n23090_o = n22438_o[42:35];
  /* mmu.vhdl:231:54  */
  assign n23091_o = n22438_o[34:27];
  /* mmu.vhdl:231:54  */
  assign n23092_o = n22438_o[26:19];
  /* mmu.vhdl:231:54  */
  assign n23093_o = n22438_o[18:11];
  /* mmu.vhdl:231:54  */
  assign n23094_o = n22438_o[10:3];
  /* mmu.vhdl:234:16  */
  assign n23095_o = r[168:165];
  /* mmu.vhdl:236:25  */
  assign n23096_o = n22421_o[80];
  /* mmu.vhdl:236:30  */
  assign n23097_o = ~n23096_o;
  /* mmu.vhdl:237:28  */
  assign n23098_o = r[299:236];
  /* mmu.vhdl:238:31  */
  assign n23099_o = r[300];
  /* mmu.vhdl:240:28  */
  assign n23100_o = r[364:301];
  /* mmu.vhdl:241:31  */
  assign n23101_o = r[365];
  /* mmu.vhdl:236:13  */
  assign n23102_o = n23097_o ? n23099_o : n23101_o;
  /* mmu.vhdl:236:13  */
  assign n23103_o = n23097_o ? n23098_o : n23100_o;
  /* mmu.vhdl:244:40  */
  assign n23104_o = n23103_o[62:61];
  /* mmu.vhdl:244:33  */
  assign n23106_o = {1'b0, n23104_o};
  /* mmu.vhdl:244:62  */
  assign n23107_o = n23103_o[7:5];
  /* mmu.vhdl:244:55  */
  assign n23108_o = {n23106_o, n23107_o};
  /* mmu.vhdl:246:42  */
  assign n23109_o = n23103_o[4:0];
  /* mmu.vhdl:246:35  */
  assign n23111_o = {1'b0, n23109_o};
  /* mmu.vhdl:249:33  */
  assign n23112_o = n23111_o[4:0];
  /* mmu.vhdl:250:30  */
  assign n23113_o = n23103_o[55:8];
  /* mmu.vhdl:250:44  */
  assign n23115_o = {n23113_o, 8'b00000000};
  /* mmu.vhdl:252:21  */
  assign n23116_o = n22421_o[0];
  /* mmu.vhdl:253:32  */
  assign n23117_o = n22421_o[80:17];
  /* mmu.vhdl:254:33  */
  assign n23118_o = n22421_o[4];
  /* mmu.vhdl:255:38  */
  assign n23119_o = n22421_o[5];
  /* mmu.vhdl:255:51  */
  assign n23120_o = n22421_o[4];
  /* mmu.vhdl:255:43  */
  assign n23121_o = n23119_o | n23120_o;
  /* mmu.vhdl:255:28  */
  assign n23122_o = ~n23121_o;
  /* mmu.vhdl:256:32  */
  assign n23123_o = n22421_o[6];
  /* mmu.vhdl:257:25  */
  assign n23124_o = n22421_o[1];
  /* mmu.vhdl:260:41  */
  assign n23125_o = n22421_o[2];
  /* mmu.vhdl:260:59  */
  assign n23126_o = n22421_o[28];
  /* mmu.vhdl:260:47  */
  assign n23127_o = n23125_o | n23126_o;
  /* mmu.vhdl:260:76  */
  assign n23128_o = n22421_o[27];
  /* mmu.vhdl:260:64  */
  assign n23129_o = n23127_o | n23128_o;
  /* mmu.vhdl:261:45  */
  assign n23130_o = n22421_o[24];
  /* mmu.vhdl:260:81  */
  assign n23131_o = n23129_o | n23130_o;
  /* mmu.vhdl:261:61  */
  assign n23132_o = n22421_o[23];
  /* mmu.vhdl:261:49  */
  assign n23133_o = n23131_o | n23132_o;
  /* mmu.vhdl:261:77  */
  assign n23134_o = n22421_o[22];
  /* mmu.vhdl:261:65  */
  assign n23135_o = n23133_o | n23134_o;
  /* mmu.vhdl:264:33  */
  assign n23136_o = n22421_o[10];
  assign n23140_o = r[235];
  /* mmu.vhdl:252:13  */
  assign n23141_o = n23187_o ? 1'b0 : n23140_o;
  assign n23142_o = r[300];
  /* mmu.vhdl:252:13  */
  assign n23143_o = n23189_o ? 1'b0 : n23142_o;
  assign n23144_o = r[365];
  /* mmu.vhdl:257:17  */
  assign n23145_o = n23177_o ? 1'b0 : n23144_o;
  /* mmu.vhdl:272:26  */
  assign n23148_o = r[235];
  /* mmu.vhdl:272:36  */
  assign n23149_o = ~n23148_o;
  /* mmu.vhdl:275:36  */
  assign n23151_o = ~n23102_o;
  /* mmu.vhdl:279:58  */
  assign n23152_o = r[175:171];
  /* mmu.vhdl:279:49  */
  assign n23154_o = {1'b0, n23152_o};
  /* mmu.vhdl:281:33  */
  assign n23157_o = n23111_o == 6'b000000;
  /* mmu.vhdl:281:21  */
  assign n23161_o = n23157_o ? 4'b1100 : 4'b1000;
  /* mmu.vhdl:281:21  */
  assign n23162_o = n23157_o ? 1'b1 : 1'b0;
  /* mmu.vhdl:275:21  */
  assign n23163_o = n23151_o ? 4'b0110 : n23161_o;
  /* mmu.vhdl:275:21  */
  assign n23164_o = n23151_o ? n23154_o : n23108_o;
  /* mmu.vhdl:275:21  */
  assign n23165_o = n23151_o ? 1'b0 : n23162_o;
  /* mmu.vhdl:272:21  */
  assign n23166_o = n23149_o ? 4'b0011 : n23163_o;
  /* mmu.vhdl:272:21  */
  assign n23167_o = n23149_o ? n23108_o : n23164_o;
  /* mmu.vhdl:272:21  */
  assign n23168_o = n23149_o ? 1'b0 : n23165_o;
  /* mmu.vhdl:257:17  */
  assign n23169_o = n23124_o ? 1'b0 : 1'b1;
  /* mmu.vhdl:257:17  */
  assign n23170_o = n23124_o ? n23135_o : 1'b0;
  /* mmu.vhdl:257:17  */
  assign n23171_o = n23124_o ? 4'b0001 : n23166_o;
  /* mmu.vhdl:257:17  */
  assign n23173_o = n23124_o & n23136_o;
  /* mmu.vhdl:257:17  */
  assign n23175_o = n23124_o & n23136_o;
  /* mmu.vhdl:257:17  */
  assign n23177_o = n23124_o & n23136_o;
  /* mmu.vhdl:257:17  */
  assign n23178_o = n23124_o ? n23108_o : n23167_o;
  /* mmu.vhdl:257:17  */
  assign n23179_o = n23124_o ? 1'b0 : n23168_o;
  assign n23180_o = {n23170_o, n23117_o, n23123_o, n23122_o, n23118_o, n23169_o};
  assign n23181_o = {n23178_o, n23145_o};
  assign n23182_o = {1'b0, n23086_o, 1'b0};
  assign n23184_o = r[168:165];
  /* mmu.vhdl:252:13  */
  assign n23185_o = n23116_o ? n23171_o : n23184_o;
  /* mmu.vhdl:252:13  */
  assign n23187_o = n23116_o & n23173_o;
  /* mmu.vhdl:252:13  */
  assign n23189_o = n23116_o & n23175_o;
  assign n23190_o = r[365];
  assign n23191_o = {n23108_o, n23190_o};
  /* mmu.vhdl:252:13  */
  assign n23193_o = n23116_o ? n23179_o : 1'b0;
  /* mmu.vhdl:290:21  */
  assign n23194_o = n22421_o[3];
  /* mmu.vhdl:294:29  */
  assign n23195_o = n22421_o[15];
  /* mmu.vhdl:294:33  */
  assign n23196_o = ~n23195_o;
  /* mmu.vhdl:295:37  */
  assign n23197_o = n22421_o[112:81];
  /* mmu.vhdl:297:36  */
  assign n23198_o = n22421_o[144:81];
  assign n23201_o = r[132:69];
  /* mmu.vhdl:294:17  */
  assign n23202_o = n23196_o ? n23201_o : n23198_o;
  assign n23203_o = r[164:133];
  /* mmu.vhdl:294:17  */
  assign n23204_o = n23196_o ? n23197_o : n23203_o;
  /* mmu.vhdl:294:17  */
  assign n23205_o = n23196_o ? n23141_o : 1'b0;
  assign n23206_o = n23181_o[0];
  assign n23207_o = n23191_o[0];
  /* mmu.vhdl:252:13  */
  assign n23208_o = n23116_o ? n23206_o : n23207_o;
  /* mmu.vhdl:294:17  */
  assign n23209_o = n23196_o ? n23208_o : 1'b0;
  assign n23213_o = {4'b0001, n23204_o, n23202_o, 1'b1};
  assign n23214_o = n23180_o[68];
  assign n23215_o = n23182_o[68];
  /* mmu.vhdl:252:13  */
  assign n23216_o = n23116_o ? n23214_o : n23215_o;
  assign n23217_o = r[164:69];
  assign n23218_o = {n23185_o, n23217_o, n23216_o};
  /* mmu.vhdl:290:13  */
  assign n23219_o = n23194_o ? n23213_o : n23218_o;
  /* mmu.vhdl:290:13  */
  assign n23220_o = n23194_o ? n23205_o : n23141_o;
  /* mmu.vhdl:290:13  */
  assign n23221_o = n23194_o ? 1'b0 : n23143_o;
  assign n23222_o = n23181_o[0];
  assign n23223_o = n23191_o[0];
  /* mmu.vhdl:252:13  */
  assign n23224_o = n23116_o ? n23222_o : n23223_o;
  /* mmu.vhdl:290:13  */
  assign n23225_o = n23194_o ? n23209_o : n23224_o;
  assign n23226_o = n23180_o[67:0];
  assign n23227_o = n23182_o[67:0];
  /* mmu.vhdl:252:13  */
  assign n23228_o = n23116_o ? n23226_o : n23227_o;
  assign n23229_o = n23181_o[6:1];
  assign n23230_o = n23191_o[6:1];
  /* mmu.vhdl:252:13  */
  assign n23231_o = n23116_o ? n23229_o : n23230_o;
  /* mmu.vhdl:235:9  */
  assign n23233_o = n23095_o == 4'b0000;
  /* mmu.vhdl:306:9  */
  assign n23236_o = n23095_o == 4'b0001;
  /* mmu.vhdl:312:21  */
  assign n23237_o = n22438_o[1];
  assign n23239_o = r[168:165];
  /* mmu.vhdl:312:13  */
  assign n23240_o = n23237_o ? 4'b1100 : n23239_o;
  /* mmu.vhdl:311:9  */
  assign n23242_o = n23095_o == 4'b0010;
  /* mmu.vhdl:316:9  */
  assign n23245_o = n23095_o == 4'b0011;
  /* mmu.vhdl:322:21  */
  assign n23246_o = n22438_o[1];
  assign n23247_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  assign n23250_o = {1'b1, n23247_o};
  assign n23251_o = r[168:165];
  /* mmu.vhdl:322:13  */
  assign n23252_o = n23246_o ? 4'b0101 : n23251_o;
  assign n23253_o = r[235:171];
  /* mmu.vhdl:322:13  */
  assign n23254_o = n23246_o ? n23250_o : n23253_o;
  /* mmu.vhdl:321:9  */
  assign n23256_o = n23095_o == 4'b0100;
  /* mmu.vhdl:329:46  */
  assign n23257_o = r[175:171];
  /* mmu.vhdl:329:37  */
  assign n23259_o = {1'b0, n23257_o};
  /* mmu.vhdl:328:9  */
  assign n23262_o = n23095_o == 4'b0101;
  /* mmu.vhdl:332:9  */
  assign n23265_o = n23095_o == 4'b0110;
  /* mmu.vhdl:338:21  */
  assign n23266_o = n22438_o[1];
  /* mmu.vhdl:339:26  */
  assign n23267_o = r[67];
  assign n23268_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  assign n23270_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  assign n23272_o = {1'b1, n23270_o};
  assign n23273_o = {1'b1, n23268_o};
  assign n23274_o = r[300:236];
  /* mmu.vhdl:339:17  */
  assign n23275_o = n23267_o ? n23274_o : n23272_o;
  assign n23276_o = r[365:301];
  /* mmu.vhdl:339:17  */
  assign n23277_o = n23267_o ? n23273_o : n23276_o;
  assign n23278_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:347:43  */
  assign n23279_o = n23278_o[62:61];
  /* mmu.vhdl:347:37  */
  assign n23281_o = {1'b0, n23279_o};
  assign n23282_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:347:64  */
  assign n23283_o = n23282_o[7:5];
  /* mmu.vhdl:347:58  */
  assign n23284_o = {n23281_o, n23283_o};
  assign n23285_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:349:45  */
  assign n23286_o = n23285_o[4:0];
  /* mmu.vhdl:349:39  */
  assign n23288_o = {1'b0, n23286_o};
  /* mmu.vhdl:352:37  */
  assign n23289_o = n23288_o[4:0];
  assign n23290_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:353:33  */
  assign n23291_o = n23290_o[55:8];
  /* mmu.vhdl:353:47  */
  assign n23293_o = {n23291_o, 8'b00000000};
  /* mmu.vhdl:354:26  */
  assign n23295_o = n23288_o == 6'b000000;
  /* mmu.vhdl:354:17  */
  assign n23299_o = n23295_o ? 4'b1100 : 4'b1000;
  /* mmu.vhdl:338:13  */
  assign n23300_o = n23306_o ? 1'b1 : 1'b0;
  assign n23301_o = {n23293_o, n23289_o, n23284_o, n23277_o, n23275_o};
  assign n23302_o = r[168:165];
  /* mmu.vhdl:338:13  */
  assign n23303_o = n23266_o ? n23299_o : n23302_o;
  assign n23304_o = r[432:236];
  /* mmu.vhdl:338:13  */
  assign n23305_o = n23266_o ? n23301_o : n23304_o;
  /* mmu.vhdl:338:13  */
  assign n23306_o = n23266_o & n23295_o;
  /* mmu.vhdl:361:21  */
  assign n23309_o = n22438_o[2];
  /* mmu.vhdl:361:13  */
  assign n23312_o = n23309_o ? 4'b1100 : n23303_o;
  /* mmu.vhdl:361:13  */
  assign n23313_o = n23309_o ? 1'b1 : 1'b0;
  /* mmu.vhdl:337:9  */
  assign n23315_o = n23095_o == 4'b0111;
  /* mmu.vhdl:367:30  */
  assign n23316_o = r[376:372];
  /* mmu.vhdl:367:26  */
  assign n23318_o = {1'b0, n23316_o};
  /* mmu.vhdl:368:26  */
  assign n23319_o = r[371:366];
  /* mmu.vhdl:368:32  */
  assign n23321_o = n23319_o + 6'b010011;
  /* mmu.vhdl:368:44  */
  assign n23322_o = n23321_o - n23318_o;
  /* mmu.vhdl:369:33  */
  assign n23323_o = r[65:35];
  /* mmu.vhdl:369:65  */
  assign n23324_o = finalmask[30:0];
  /* mmu.vhdl:369:52  */
  assign n23325_o = ~n23324_o;
  /* mmu.vhdl:369:48  */
  assign n23326_o = n23323_o & n23325_o;
  /* mmu.vhdl:369:24  */
  assign n23327_o = |(n23326_o);
  /* mmu.vhdl:370:22  */
  assign n23328_o = r[67];
  /* mmu.vhdl:370:36  */
  assign n23329_o = r[66];
  /* mmu.vhdl:370:27  */
  assign n23330_o = n23328_o != n23329_o;
  /* mmu.vhdl:370:41  */
  assign n23331_o = n23330_o | n23327_o;
  /* mmu.vhdl:373:25  */
  assign n23335_o = $unsigned(n23318_o) < $unsigned(6'b000101);
  /* mmu.vhdl:373:38  */
  assign n23337_o = $unsigned(n23318_o) > $unsigned(6'b010000);
  /* mmu.vhdl:373:29  */
  assign n23338_o = n23335_o | n23337_o;
  /* mmu.vhdl:373:57  */
  assign n23339_o = r[371:366];
  /* mmu.vhdl:373:63  */
  assign n23341_o = n23339_o + 6'b010011;
  /* mmu.vhdl:373:52  */
  assign n23342_o = $unsigned(n23318_o) > $unsigned(n23341_o);
  /* mmu.vhdl:373:43  */
  assign n23343_o = n23338_o | n23342_o;
  /* mmu.vhdl:373:13  */
  assign n23347_o = n23343_o ? 4'b1100 : 4'b1001;
  /* mmu.vhdl:373:13  */
  assign n23348_o = n23343_o ? 1'b1 : 1'b0;
  /* mmu.vhdl:370:13  */
  assign n23349_o = n23331_o ? 4'b1100 : n23347_o;
  /* mmu.vhdl:370:13  */
  assign n23350_o = n23331_o ? 1'b0 : n23348_o;
  /* mmu.vhdl:370:13  */
  assign n23351_o = n23331_o ? 1'b1 : 1'b0;
  /* mmu.vhdl:366:9  */
  assign n23353_o = n23095_o == 4'b1000;
  /* mmu.vhdl:380:9  */
  assign n23356_o = n23095_o == 4'b1001;
  /* mmu.vhdl:385:21  */
  assign n23357_o = n22438_o[1];
  assign n23358_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  assign n23359_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:388:24  */
  assign n23360_o = n23359_o[63];
  assign n23361_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:390:28  */
  assign n23362_o = n23361_o[62];
  /* mmu.vhdl:393:30  */
  assign n23363_o = r[3];
  assign n23364_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:393:48  */
  assign n23365_o = n23364_o[3];
  /* mmu.vhdl:393:52  */
  assign n23366_o = ~n23365_o;
  /* mmu.vhdl:393:41  */
  assign n23367_o = n23363_o | n23366_o;
  /* mmu.vhdl:394:34  */
  assign n23368_o = r[1];
  /* mmu.vhdl:394:40  */
  assign n23369_o = ~n23368_o;
  assign n23370_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:395:48  */
  assign n23371_o = n23370_o[1];
  assign n23372_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:395:60  */
  assign n23373_o = n23372_o[2];
  /* mmu.vhdl:395:74  */
  assign n23374_o = r[2];
  /* mmu.vhdl:395:68  */
  assign n23375_o = ~n23374_o;
  /* mmu.vhdl:395:64  */
  assign n23376_o = n23373_o & n23375_o;
  /* mmu.vhdl:395:52  */
  assign n23377_o = n23371_o | n23376_o;
  assign n23378_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:399:48  */
  assign n23379_o = n23378_o[0];
  assign n23380_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:399:64  */
  assign n23381_o = n23380_o[5];
  /* mmu.vhdl:399:56  */
  assign n23382_o = ~n23381_o;
  /* mmu.vhdl:399:52  */
  assign n23383_o = n23379_o & n23382_o;
  /* mmu.vhdl:394:29  */
  assign n23384_o = n23369_o ? n23377_o : n23383_o;
  /* mmu.vhdl:393:25  */
  assign n23386_o = n23367_o ? n23384_o : 1'b0;
  assign n23388_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:402:38  */
  assign n23389_o = n23388_o[8];
  assign n23390_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:402:51  */
  assign n23391_o = n23390_o[7];
  /* mmu.vhdl:402:64  */
  assign n23392_o = r[2];
  /* mmu.vhdl:402:58  */
  assign n23393_o = ~n23392_o;
  /* mmu.vhdl:402:55  */
  assign n23394_o = n23391_o | n23393_o;
  /* mmu.vhdl:402:42  */
  assign n23395_o = n23389_o & n23394_o;
  /* mmu.vhdl:403:42  */
  assign n23396_o = n23386_o & n23395_o;
  /* mmu.vhdl:407:43  */
  assign n23399_o = ~n23386_o;
  assign n23400_o = {n23386_o, n23399_o};
  /* mmu.vhdl:403:25  */
  assign n23401_o = n23396_o ? 4'b1011 : 4'b1100;
  assign n23402_o = {1'b0, 1'b0};
  /* mmu.vhdl:403:25  */
  assign n23403_o = n23396_o ? n23402_o : n23400_o;
  assign n23404_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:412:53  */
  assign n23405_o = n23404_o[4:0];
  /* mmu.vhdl:412:47  */
  assign n23407_o = {1'b0, n23405_o};
  /* mmu.vhdl:413:34  */
  assign n23409_o = $unsigned(n23407_o) < $unsigned(6'b000101);
  /* mmu.vhdl:413:47  */
  assign n23411_o = $unsigned(n23407_o) > $unsigned(6'b010000);
  /* mmu.vhdl:413:38  */
  assign n23412_o = n23409_o | n23411_o;
  /* mmu.vhdl:413:65  */
  assign n23413_o = r[371:366];
  /* mmu.vhdl:413:61  */
  assign n23414_o = $unsigned(n23407_o) > $unsigned(n23413_o);
  /* mmu.vhdl:413:52  */
  assign n23415_o = n23412_o | n23414_o;
  assign n23418_o = r[432:171];
  assign n23419_o = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n23358_o, n23418_o, 1'b0, 1'b0, n23085_o, 1'b0, n23086_o, 1'b0};
  /* mmu.vhdl:417:42  */
  assign n23420_o = n23419_o[371:366];
  /* mmu.vhdl:417:48  */
  assign n23421_o = n23420_o - n23407_o;
  /* mmu.vhdl:418:49  */
  assign n23422_o = n23407_o[4:0];
  assign n23423_o = {n23094_o, n23093_o, n23092_o, n23091_o, n23090_o, n23089_o, n23088_o, n23087_o};
  /* mmu.vhdl:419:45  */
  assign n23424_o = n23423_o[55:8];
  /* mmu.vhdl:419:59  */
  assign n23426_o = {n23424_o, 8'b00000000};
  assign n23428_o = {n23426_o, n23422_o, n23421_o};
  /* mmu.vhdl:413:25  */
  assign n23429_o = n23415_o ? 4'b1100 : 4'b1001;
  assign n23430_o = r[432:366];
  /* mmu.vhdl:413:25  */
  assign n23431_o = n23415_o ? n23430_o : n23428_o;
  /* mmu.vhdl:413:25  */
  assign n23432_o = n23415_o ? 1'b1 : 1'b0;
  /* mmu.vhdl:390:21  */
  assign n23433_o = n23362_o ? n23401_o : n23429_o;
  assign n23434_o = r[432:366];
  /* mmu.vhdl:390:21  */
  assign n23435_o = n23362_o ? n23434_o : n23431_o;
  /* mmu.vhdl:390:21  */
  assign n23436_o = n23362_o ? 1'b0 : n23432_o;
  assign n23437_o = {1'b0, 1'b0};
  /* mmu.vhdl:390:21  */
  assign n23438_o = n23362_o ? n23403_o : n23437_o;
  /* mmu.vhdl:388:17  */
  assign n23444_o = n23360_o ? n23433_o : 4'b1100;
  assign n23445_o = r[432:366];
  /* mmu.vhdl:388:17  */
  assign n23446_o = n23360_o ? n23435_o : n23445_o;
  /* mmu.vhdl:388:17  */
  assign n23447_o = n23360_o ? 1'b0 : 1'b1;
  /* mmu.vhdl:388:17  */
  assign n23448_o = n23360_o ? n23436_o : 1'b0;
  assign n23449_o = {1'b0, 1'b0};
  /* mmu.vhdl:388:17  */
  assign n23450_o = n23360_o ? n23438_o : n23449_o;
  assign n23454_o = {n23448_o, n23447_o, n23358_o, n23446_o};
  assign n23455_o = r[168:165];
  /* mmu.vhdl:385:13  */
  assign n23456_o = n23357_o ? n23444_o : n23455_o;
  assign n23457_o = r[496:366];
  assign n23458_o = {1'b0, 1'b0, n23457_o};
  assign n23460_o = {1'b0, 1'b0};
  /* mmu.vhdl:385:13  */
  assign n23461_o = n23357_o ? n23450_o : n23460_o;
  /* mmu.vhdl:429:21  */
  assign n23465_o = n22438_o[2];
  /* mmu.vhdl:429:13  */
  assign n23468_o = n23465_o ? 4'b1100 : n23456_o;
  assign n23469_o = n23454_o[132];
  assign n23470_o = n23458_o[132];
  /* mmu.vhdl:385:13  */
  assign n23471_o = n23357_o ? n23469_o : n23470_o;
  /* mmu.vhdl:429:13  */
  assign n23472_o = n23465_o ? 1'b1 : n23471_o;
  assign n23473_o = n23454_o[131:0];
  assign n23474_o = n23458_o[131:0];
  /* mmu.vhdl:385:13  */
  assign n23475_o = n23357_o ? n23473_o : n23474_o;
  /* mmu.vhdl:384:9  */
  assign n23477_o = n23095_o == 4'b1010;
  /* mmu.vhdl:436:18  */
  assign n23478_o = r[1];
  /* mmu.vhdl:436:24  */
  assign n23479_o = ~n23478_o;
  /* mmu.vhdl:436:13  */
  assign n23482_o = n23479_o ? 4'b0010 : 4'b0000;
  /* mmu.vhdl:436:13  */
  assign n23485_o = n23479_o ? 1'b1 : 1'b0;
  /* mmu.vhdl:436:13  */
  assign n23488_o = n23479_o ? 1'b0 : 1'b1;
  /* mmu.vhdl:434:9  */
  assign n23490_o = n23095_o == 4'b1011;
  /* mmu.vhdl:444:9  */
  assign n23493_o = n23095_o == 4'b1100;
  assign n23494_o = {n23493_o, n23490_o, n23477_o, n23356_o, n23353_o, n23315_o, n23265_o, n23262_o, n23256_o, n23245_o, n23242_o, n23236_o, n23233_o};
  assign n23495_o = {n23086_o, 1'b0};
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23497_o = n23495_o;
      13'b0100000000000: n23497_o = n23495_o;
      13'b0010000000000: n23497_o = n23495_o;
      13'b0001000000000: n23497_o = n23495_o;
      13'b0000100000000: n23497_o = n23495_o;
      13'b0000010000000: n23497_o = n23495_o;
      13'b0000001000000: n23497_o = n23495_o;
      13'b0000000100000: n23497_o = n23495_o;
      13'b0000000010000: n23497_o = n23495_o;
      13'b0000000001000: n23497_o = n23495_o;
      13'b0000000000100: n23497_o = n23495_o;
      13'b0000000000010: n23497_o = n23495_o;
      13'b0000000000001: n23497_o = n23228_o;
      default: n23497_o = 68'bX;
    endcase
  assign n23498_o = n23219_o[96:0];
  assign n23499_o = r[164:69];
  assign n23500_o = {n23499_o, 1'b0};
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23502_o = n23500_o;
      13'b0100000000000: n23502_o = n23500_o;
      13'b0010000000000: n23502_o = n23500_o;
      13'b0001000000000: n23502_o = n23500_o;
      13'b0000100000000: n23502_o = n23500_o;
      13'b0000010000000: n23502_o = n23500_o;
      13'b0000001000000: n23502_o = n23500_o;
      13'b0000000100000: n23502_o = n23500_o;
      13'b0000000010000: n23502_o = n23500_o;
      13'b0000000001000: n23502_o = n23500_o;
      13'b0000000000100: n23502_o = n23500_o;
      13'b0000000000010: n23502_o = n23500_o;
      13'b0000000000001: n23502_o = n23498_o;
      default: n23502_o = 97'bX;
    endcase
  assign n23503_o = n23219_o[100:97];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23505_o = 4'b0000;
      13'b0100000000000: n23505_o = n23482_o;
      13'b0010000000000: n23505_o = n23468_o;
      13'b0001000000000: n23505_o = 4'b1010;
      13'b0000100000000: n23505_o = n23349_o;
      13'b0000010000000: n23505_o = n23312_o;
      13'b0000001000000: n23505_o = 4'b0111;
      13'b0000000100000: n23505_o = 4'b0110;
      13'b0000000010000: n23505_o = n23252_o;
      13'b0000000001000: n23505_o = 4'b0100;
      13'b0000000000100: n23505_o = n23240_o;
      13'b0000000000010: n23505_o = 4'b0010;
      13'b0000000000001: n23505_o = n23503_o;
      default: n23505_o = 4'bX;
    endcase
  assign n23506_o = n23254_o[63:0];
  assign n23507_o = r[234:171];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23509_o = n23507_o;
      13'b0100000000000: n23509_o = n23507_o;
      13'b0010000000000: n23509_o = n23507_o;
      13'b0001000000000: n23509_o = n23507_o;
      13'b0000100000000: n23509_o = n23507_o;
      13'b0000010000000: n23509_o = n23507_o;
      13'b0000001000000: n23509_o = n23507_o;
      13'b0000000100000: n23509_o = n23507_o;
      13'b0000000010000: n23509_o = n23506_o;
      13'b0000000001000: n23509_o = n23507_o;
      13'b0000000000100: n23509_o = n23507_o;
      13'b0000000000010: n23509_o = n23507_o;
      13'b0000000000001: n23509_o = n23507_o;
      default: n23509_o = 64'bX;
    endcase
  assign n23510_o = n23254_o[64];
  assign n23511_o = r[235];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23513_o = n23511_o;
      13'b0100000000000: n23513_o = n23511_o;
      13'b0010000000000: n23513_o = n23511_o;
      13'b0001000000000: n23513_o = n23511_o;
      13'b0000100000000: n23513_o = n23511_o;
      13'b0000010000000: n23513_o = n23511_o;
      13'b0000001000000: n23513_o = n23511_o;
      13'b0000000100000: n23513_o = n23511_o;
      13'b0000000010000: n23513_o = n23510_o;
      13'b0000000001000: n23513_o = n23511_o;
      13'b0000000000100: n23513_o = n23511_o;
      13'b0000000000010: n23513_o = n23511_o;
      13'b0000000000001: n23513_o = n23220_o;
      default: n23513_o = 1'bX;
    endcase
  assign n23514_o = n23305_o[63:0];
  assign n23515_o = r[299:236];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23517_o = n23515_o;
      13'b0100000000000: n23517_o = n23515_o;
      13'b0010000000000: n23517_o = n23515_o;
      13'b0001000000000: n23517_o = n23515_o;
      13'b0000100000000: n23517_o = n23515_o;
      13'b0000010000000: n23517_o = n23514_o;
      13'b0000001000000: n23517_o = n23515_o;
      13'b0000000100000: n23517_o = n23515_o;
      13'b0000000010000: n23517_o = n23515_o;
      13'b0000000001000: n23517_o = n23515_o;
      13'b0000000000100: n23517_o = n23515_o;
      13'b0000000000010: n23517_o = n23515_o;
      13'b0000000000001: n23517_o = n23515_o;
      default: n23517_o = 64'bX;
    endcase
  assign n23518_o = n23305_o[64];
  assign n23519_o = r[300];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23521_o = n23519_o;
      13'b0100000000000: n23521_o = n23519_o;
      13'b0010000000000: n23521_o = n23519_o;
      13'b0001000000000: n23521_o = n23519_o;
      13'b0000100000000: n23521_o = n23519_o;
      13'b0000010000000: n23521_o = n23518_o;
      13'b0000001000000: n23521_o = n23519_o;
      13'b0000000100000: n23521_o = n23519_o;
      13'b0000000010000: n23521_o = n23519_o;
      13'b0000000001000: n23521_o = n23519_o;
      13'b0000000000100: n23521_o = n23519_o;
      13'b0000000000010: n23521_o = n23519_o;
      13'b0000000000001: n23521_o = n23221_o;
      default: n23521_o = 1'bX;
    endcase
  assign n23522_o = n23305_o[128:65];
  assign n23523_o = r[364:301];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23525_o = n23523_o;
      13'b0100000000000: n23525_o = n23523_o;
      13'b0010000000000: n23525_o = n23523_o;
      13'b0001000000000: n23525_o = n23523_o;
      13'b0000100000000: n23525_o = n23523_o;
      13'b0000010000000: n23525_o = n23522_o;
      13'b0000001000000: n23525_o = n23523_o;
      13'b0000000100000: n23525_o = n23523_o;
      13'b0000000010000: n23525_o = n23523_o;
      13'b0000000001000: n23525_o = n23523_o;
      13'b0000000000100: n23525_o = n23523_o;
      13'b0000000000010: n23525_o = n23523_o;
      13'b0000000000001: n23525_o = n23523_o;
      default: n23525_o = 64'bX;
    endcase
  assign n23526_o = n23305_o[129];
  assign n23527_o = r[365];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23529_o = n23527_o;
      13'b0100000000000: n23529_o = n23527_o;
      13'b0010000000000: n23529_o = n23527_o;
      13'b0001000000000: n23529_o = n23527_o;
      13'b0000100000000: n23529_o = n23527_o;
      13'b0000010000000: n23529_o = n23526_o;
      13'b0000001000000: n23529_o = n23527_o;
      13'b0000000100000: n23529_o = n23527_o;
      13'b0000000010000: n23529_o = n23527_o;
      13'b0000000001000: n23529_o = n23527_o;
      13'b0000000000100: n23529_o = n23527_o;
      13'b0000000000010: n23529_o = n23527_o;
      13'b0000000000001: n23529_o = n23225_o;
      default: n23529_o = 1'bX;
    endcase
  assign n23530_o = n23305_o[135:130];
  assign n23531_o = n23475_o[5:0];
  assign n23532_o = r[371:366];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23534_o = n23532_o;
      13'b0100000000000: n23534_o = n23532_o;
      13'b0010000000000: n23534_o = n23531_o;
      13'b0001000000000: n23534_o = n23532_o;
      13'b0000100000000: n23534_o = n23322_o;
      13'b0000010000000: n23534_o = n23530_o;
      13'b0000001000000: n23534_o = n23532_o;
      13'b0000000100000: n23534_o = n23259_o;
      13'b0000000010000: n23534_o = n23532_o;
      13'b0000000001000: n23534_o = n23532_o;
      13'b0000000000100: n23534_o = n23532_o;
      13'b0000000000010: n23534_o = n23532_o;
      13'b0000000000001: n23534_o = n23231_o;
      default: n23534_o = 6'bX;
    endcase
  assign n23535_o = n23305_o[140:136];
  assign n23536_o = n23475_o[10:6];
  assign n23537_o = r[376:372];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23539_o = n23537_o;
      13'b0100000000000: n23539_o = n23537_o;
      13'b0010000000000: n23539_o = n23536_o;
      13'b0001000000000: n23539_o = n23537_o;
      13'b0000100000000: n23539_o = n23537_o;
      13'b0000010000000: n23539_o = n23535_o;
      13'b0000001000000: n23539_o = n23537_o;
      13'b0000000100000: n23539_o = n23537_o;
      13'b0000000010000: n23539_o = n23537_o;
      13'b0000000001000: n23539_o = n23537_o;
      13'b0000000000100: n23539_o = n23537_o;
      13'b0000000000010: n23539_o = n23537_o;
      13'b0000000000001: n23539_o = n23112_o;
      default: n23539_o = 5'bX;
    endcase
  assign n23540_o = n23305_o[196:141];
  assign n23541_o = n23475_o[66:11];
  assign n23542_o = r[432:377];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23544_o = n23542_o;
      13'b0100000000000: n23544_o = n23542_o;
      13'b0010000000000: n23544_o = n23541_o;
      13'b0001000000000: n23544_o = n23542_o;
      13'b0000100000000: n23544_o = n23542_o;
      13'b0000010000000: n23544_o = n23540_o;
      13'b0000001000000: n23544_o = n23542_o;
      13'b0000000100000: n23544_o = n23542_o;
      13'b0000000010000: n23544_o = n23542_o;
      13'b0000000001000: n23544_o = n23542_o;
      13'b0000000000100: n23544_o = n23542_o;
      13'b0000000000010: n23544_o = n23542_o;
      13'b0000000000001: n23544_o = n23115_o;
      default: n23544_o = 56'bX;
    endcase
  assign n23545_o = n23475_o[130:67];
  assign n23546_o = r[496:433];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23548_o = n23546_o;
      13'b0100000000000: n23548_o = n23546_o;
      13'b0010000000000: n23548_o = n23545_o;
      13'b0001000000000: n23548_o = n23546_o;
      13'b0000100000000: n23548_o = n23546_o;
      13'b0000010000000: n23548_o = n23546_o;
      13'b0000001000000: n23548_o = n23546_o;
      13'b0000000100000: n23548_o = n23546_o;
      13'b0000000010000: n23548_o = n23546_o;
      13'b0000000001000: n23548_o = n23546_o;
      13'b0000000000100: n23548_o = n23546_o;
      13'b0000000000010: n23548_o = n23546_o;
      13'b0000000000001: n23548_o = n23546_o;
      default: n23548_o = 64'bX;
    endcase
  assign n23549_o = n23475_o[131];
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23551_o = 1'b0;
      13'b0100000000000: n23551_o = 1'b0;
      13'b0010000000000: n23551_o = n23549_o;
      13'b0001000000000: n23551_o = 1'b0;
      13'b0000100000000: n23551_o = 1'b0;
      13'b0000010000000: n23551_o = n23300_o;
      13'b0000001000000: n23551_o = 1'b0;
      13'b0000000100000: n23551_o = 1'b0;
      13'b0000000010000: n23551_o = 1'b0;
      13'b0000000001000: n23551_o = 1'b0;
      13'b0000000000100: n23551_o = 1'b0;
      13'b0000000000010: n23551_o = 1'b0;
      13'b0000000000001: n23551_o = n23193_o;
      default: n23551_o = 1'bX;
    endcase
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23553_o = 1'b0;
      13'b0100000000000: n23553_o = 1'b0;
      13'b0010000000000: n23553_o = n23472_o;
      13'b0001000000000: n23553_o = 1'b0;
      13'b0000100000000: n23553_o = n23350_o;
      13'b0000010000000: n23553_o = n23313_o;
      13'b0000001000000: n23553_o = 1'b0;
      13'b0000000100000: n23553_o = 1'b0;
      13'b0000000010000: n23553_o = 1'b0;
      13'b0000000001000: n23553_o = 1'b0;
      13'b0000000000100: n23553_o = 1'b0;
      13'b0000000000010: n23553_o = 1'b0;
      13'b0000000000001: n23553_o = 1'b0;
      default: n23553_o = 1'bX;
    endcase
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23555_o = 1'b0;
      13'b0100000000000: n23555_o = 1'b0;
      13'b0010000000000: n23555_o = 1'b0;
      13'b0001000000000: n23555_o = 1'b0;
      13'b0000100000000: n23555_o = n23351_o;
      13'b0000010000000: n23555_o = 1'b0;
      13'b0000001000000: n23555_o = 1'b0;
      13'b0000000100000: n23555_o = 1'b0;
      13'b0000000010000: n23555_o = 1'b0;
      13'b0000000001000: n23555_o = 1'b0;
      13'b0000000000100: n23555_o = 1'b0;
      13'b0000000000010: n23555_o = 1'b0;
      13'b0000000000001: n23555_o = 1'b0;
      default: n23555_o = 1'bX;
    endcase
  assign n23556_o = {1'b0, 1'b0};
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23558_o = n23556_o;
      13'b0100000000000: n23558_o = n23556_o;
      13'b0010000000000: n23558_o = n23461_o;
      13'b0001000000000: n23558_o = n23556_o;
      13'b0000100000000: n23558_o = n23556_o;
      13'b0000010000000: n23558_o = n23556_o;
      13'b0000001000000: n23558_o = n23556_o;
      13'b0000000100000: n23558_o = n23556_o;
      13'b0000000010000: n23558_o = n23556_o;
      13'b0000000001000: n23558_o = n23556_o;
      13'b0000000000100: n23558_o = n23556_o;
      13'b0000000000010: n23558_o = n23556_o;
      13'b0000000000001: n23558_o = n23556_o;
      default: n23558_o = 2'bX;
    endcase
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23575_o = 1'b0;
      13'b0100000000000: n23575_o = n23485_o;
      13'b0010000000000: n23575_o = 1'b0;
      13'b0001000000000: n23575_o = 1'b1;
      13'b0000100000000: n23575_o = 1'b0;
      13'b0000010000000: n23575_o = 1'b0;
      13'b0000001000000: n23575_o = 1'b1;
      13'b0000000100000: n23575_o = 1'b0;
      13'b0000000010000: n23575_o = 1'b0;
      13'b0000000001000: n23575_o = 1'b1;
      13'b0000000000100: n23575_o = 1'b0;
      13'b0000000000010: n23575_o = 1'b1;
      13'b0000000000001: n23575_o = 1'b0;
      default: n23575_o = 1'bX;
    endcase
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23580_o = 1'b0;
      13'b0100000000000: n23580_o = 1'b1;
      13'b0010000000000: n23580_o = 1'b0;
      13'b0001000000000: n23580_o = 1'b0;
      13'b0000100000000: n23580_o = 1'b0;
      13'b0000010000000: n23580_o = 1'b0;
      13'b0000001000000: n23580_o = 1'b0;
      13'b0000000100000: n23580_o = 1'b0;
      13'b0000000010000: n23580_o = 1'b0;
      13'b0000000001000: n23580_o = 1'b0;
      13'b0000000000100: n23580_o = 1'b0;
      13'b0000000000010: n23580_o = 1'b0;
      13'b0000000000001: n23580_o = 1'b0;
      default: n23580_o = 1'bX;
    endcase
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23584_o = 1'b0;
      13'b0100000000000: n23584_o = n23488_o;
      13'b0010000000000: n23584_o = 1'b0;
      13'b0001000000000: n23584_o = 1'b0;
      13'b0000100000000: n23584_o = 1'b0;
      13'b0000010000000: n23584_o = 1'b0;
      13'b0000001000000: n23584_o = 1'b0;
      13'b0000000100000: n23584_o = 1'b0;
      13'b0000000010000: n23584_o = 1'b0;
      13'b0000000001000: n23584_o = 1'b0;
      13'b0000000000100: n23584_o = 1'b0;
      13'b0000000000010: n23584_o = 1'b0;
      13'b0000000000001: n23584_o = 1'b0;
      default: n23584_o = 1'bX;
    endcase
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23589_o = 1'b0;
      13'b0100000000000: n23589_o = 1'b0;
      13'b0010000000000: n23589_o = 1'b0;
      13'b0001000000000: n23589_o = 1'b0;
      13'b0000100000000: n23589_o = 1'b0;
      13'b0000010000000: n23589_o = 1'b0;
      13'b0000001000000: n23589_o = 1'b0;
      13'b0000000100000: n23589_o = 1'b0;
      13'b0000000010000: n23589_o = 1'b0;
      13'b0000000001000: n23589_o = 1'b0;
      13'b0000000000100: n23589_o = 1'b0;
      13'b0000000000010: n23589_o = 1'b1;
      13'b0000000000001: n23589_o = 1'b0;
      default: n23589_o = 1'bX;
    endcase
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23594_o = 1'b0;
      13'b0100000000000: n23594_o = 1'b0;
      13'b0010000000000: n23594_o = 1'b0;
      13'b0001000000000: n23594_o = 1'b0;
      13'b0000100000000: n23594_o = 1'b0;
      13'b0000010000000: n23594_o = 1'b0;
      13'b0000001000000: n23594_o = 1'b0;
      13'b0000000100000: n23594_o = 1'b0;
      13'b0000000010000: n23594_o = 1'b0;
      13'b0000000001000: n23594_o = 1'b1;
      13'b0000000000100: n23594_o = 1'b0;
      13'b0000000000010: n23594_o = 1'b0;
      13'b0000000000001: n23594_o = 1'b0;
      default: n23594_o = 1'bX;
    endcase
  /* mmu.vhdl:234:9  */
  always @*
    case (n23494_o)
      13'b1000000000000: n23599_o = 1'b0;
      13'b0100000000000: n23599_o = 1'b0;
      13'b0010000000000: n23599_o = 1'b0;
      13'b0001000000000: n23599_o = 1'b0;
      13'b0000100000000: n23599_o = 1'b0;
      13'b0000010000000: n23599_o = 1'b0;
      13'b0000001000000: n23599_o = 1'b1;
      13'b0000000100000: n23599_o = 1'b0;
      13'b0000000010000: n23599_o = 1'b0;
      13'b0000000001000: n23599_o = 1'b0;
      13'b0000000000100: n23599_o = 1'b0;
      13'b0000000000010: n23599_o = 1'b0;
      13'b0000000000001: n23599_o = 1'b0;
      default: n23599_o = 1'bX;
    endcase
  assign n23615_o = {n23558_o, n23555_o, n23553_o, n23551_o, n23548_o, n23544_o, n23539_o, n23534_o, n23529_o, n23525_o, n23521_o, n23517_o, n23513_o, n23509_o, 1'b0, 1'b0, n23505_o, n23502_o, n23497_o};
  /* mmu.vhdl:449:14  */
  assign n23616_o = n23615_o[168:165];
  /* mmu.vhdl:449:20  */
  assign n23618_o = n23616_o == 4'b1100;
  assign n23619_o = {n23558_o, n23555_o, n23553_o, n23551_o, n23548_o, n23544_o, n23539_o, n23534_o, n23529_o, n23525_o, n23521_o, n23517_o, n23513_o, n23509_o, 1'b0, 1'b0, n23505_o, n23502_o, n23497_o};
  /* mmu.vhdl:449:41  */
  assign n23620_o = n23619_o[168:165];
  /* mmu.vhdl:449:47  */
  assign n23622_o = n23620_o == 4'b1011;
  /* mmu.vhdl:449:70  */
  assign n23623_o = r[1];
  /* mmu.vhdl:449:64  */
  assign n23624_o = n23622_o & n23623_o;
  /* mmu.vhdl:449:35  */
  assign n23625_o = n23618_o | n23624_o;
  assign n23626_o = {n23558_o, n23555_o, n23553_o, n23551_o, n23548_o, n23544_o, n23539_o, n23534_o, n23529_o, n23525_o, n23521_o, n23517_o, n23513_o, n23509_o, 1'b0, 1'b0, n23505_o, n23502_o, n23497_o};
  /* mmu.vhdl:450:24  */
  assign n23627_o = n23626_o[497];
  assign n23628_o = {n23558_o, n23555_o, n23553_o, n23551_o, n23548_o, n23544_o, n23539_o, n23534_o, n23529_o, n23525_o, n23521_o, n23517_o, n23513_o, n23509_o, 1'b0, 1'b0, n23505_o, n23502_o, n23497_o};
  /* mmu.vhdl:450:37  */
  assign n23629_o = n23628_o[498];
  /* mmu.vhdl:450:32  */
  assign n23630_o = n23627_o | n23629_o;
  assign n23631_o = {n23558_o, n23555_o, n23553_o, n23551_o, n23548_o, n23544_o, n23539_o, n23534_o, n23529_o, n23525_o, n23521_o, n23517_o, n23513_o, n23509_o, 1'b0, 1'b0, n23505_o, n23502_o, n23497_o};
  /* mmu.vhdl:450:50  */
  assign n23632_o = n23631_o[499];
  /* mmu.vhdl:450:45  */
  assign n23633_o = n23630_o | n23632_o;
  assign n23634_o = {n23558_o, n23555_o, n23553_o, n23551_o, n23548_o, n23544_o, n23539_o, n23534_o, n23529_o, n23525_o, n23521_o, n23517_o, n23513_o, n23509_o, 1'b0, 1'b0, n23505_o, n23502_o, n23497_o};
  /* mmu.vhdl:450:64  */
  assign n23635_o = n23634_o[500];
  /* mmu.vhdl:450:59  */
  assign n23636_o = n23633_o | n23635_o;
  assign n23637_o = {n23558_o, n23555_o, n23553_o, n23551_o, n23548_o, n23544_o, n23539_o, n23534_o, n23529_o, n23525_o, n23521_o, n23517_o, n23513_o, n23509_o, 1'b0, 1'b0, n23505_o, n23502_o, n23497_o};
  /* mmu.vhdl:450:78  */
  assign n23638_o = n23637_o[501];
  /* mmu.vhdl:450:73  */
  assign n23639_o = n23636_o | n23638_o;
  assign n23640_o = {n23558_o, n23555_o, n23553_o, n23551_o, n23548_o, n23544_o, n23539_o, n23534_o, n23529_o, n23525_o, n23521_o, n23517_o, n23513_o, n23509_o, n23639_o, 1'b0, n23505_o, n23502_o, n23497_o};
  /* mmu.vhdl:451:29  */
  assign n23641_o = n23640_o[170];
  /* mmu.vhdl:451:23  */
  assign n23642_o = ~n23641_o;
  assign n23643_o = {n23639_o, n23642_o};
  assign n23644_o = {1'b0, 1'b0};
  /* mmu.vhdl:449:9  */
  assign n23645_o = n23625_o ? n23643_o : n23644_o;
  /* mmu.vhdl:454:18  */
  assign n23646_o = r[67];
  /* mmu.vhdl:457:25  */
  assign n23647_o = r[164:133];
  /* mmu.vhdl:454:9  */
  assign n23649_o = n23646_o ? 32'b00000000000000000000000000000000 : n23647_o;
  /* mmu.vhdl:459:40  */
  assign n23650_o = r[226:207];
  /* mmu.vhdl:459:31  */
  assign n23652_o = {8'b00000000, n23650_o};
  /* mmu.vhdl:460:34  */
  assign n23653_o = r[206:183];
  /* mmu.vhdl:460:66  */
  assign n23654_o = finalmask[23:0];
  /* mmu.vhdl:460:53  */
  assign n23655_o = ~n23654_o;
  /* mmu.vhdl:460:49  */
  assign n23656_o = n23653_o & n23655_o;
  /* mmu.vhdl:461:33  */
  assign n23657_o = n23649_o[31:8];
  /* mmu.vhdl:461:60  */
  assign n23658_o = finalmask[23:0];
  /* mmu.vhdl:461:47  */
  assign n23659_o = n23657_o & n23658_o;
  /* mmu.vhdl:460:81  */
  assign n23660_o = n23656_o | n23659_o;
  /* mmu.vhdl:459:55  */
  assign n23661_o = {n23652_o, n23660_o};
  /* mmu.vhdl:462:31  */
  assign n23662_o = n23649_o[7:0];
  /* mmu.vhdl:461:76  */
  assign n23663_o = {n23661_o, n23662_o};
  /* mmu.vhdl:462:44  */
  assign n23665_o = {n23663_o, 4'b0000};
  /* mmu.vhdl:464:41  */
  assign n23666_o = r[432:396];
  /* mmu.vhdl:464:31  */
  assign n23668_o = {8'b00000000, n23666_o};
  /* mmu.vhdl:465:35  */
  assign n23669_o = r[395:380];
  /* mmu.vhdl:465:53  */
  assign n23670_o = ~mask;
  /* mmu.vhdl:465:49  */
  assign n23671_o = n23669_o & n23670_o;
  /* mmu.vhdl:465:74  */
  assign n23672_o = addrsh & mask;
  /* mmu.vhdl:465:63  */
  assign n23673_o = n23671_o | n23672_o;
  /* mmu.vhdl:464:56  */
  assign n23674_o = {n23668_o, n23673_o};
  /* mmu.vhdl:465:85  */
  assign n23676_o = {n23674_o, 3'b000};
  /* mmu.vhdl:468:23  */
  assign n23677_o = r[488:445];
  /* mmu.vhdl:468:42  */
  assign n23678_o = ~finalmask;
  /* mmu.vhdl:468:38  */
  assign n23679_o = n23677_o & n23678_o;
  /* mmu.vhdl:468:67  */
  assign n23680_o = r[59:16];
  /* mmu.vhdl:468:82  */
  assign n23681_o = n23680_o & finalmask;
  /* mmu.vhdl:468:57  */
  assign n23682_o = n23679_o | n23681_o;
  /* mmu.vhdl:467:22  */
  assign n23684_o = {8'b00000000, n23682_o};
  /* mmu.vhdl:469:23  */
  assign n23685_o = r[444:433];
  /* mmu.vhdl:469:16  */
  assign n23686_o = {n23684_o, n23685_o};
  assign n23687_o = {n23558_o, n23555_o, n23553_o, n23551_o, n23548_o, n23544_o, n23539_o, n23534_o, n23529_o, n23525_o, n23521_o, n23517_o, n23513_o, n23509_o, n23645_o, n23505_o, n23502_o, n23497_o};
  /* mmu.vhdl:476:23  */
  assign n23688_o = r[67:4];
  /* mmu.vhdl:479:27  */
  assign n23689_o = r[67:16];
  /* mmu.vhdl:479:42  */
  assign n23691_o = {n23689_o, 12'b000000000000};
  /* mmu.vhdl:482:35  */
  assign n23692_o = r[124:81];
  /* mmu.vhdl:482:27  */
  assign n23694_o = {8'b00000000, n23692_o};
  /* mmu.vhdl:482:50  */
  assign n23696_o = {n23694_o, 12'b000000001000};
  /* mmu.vhdl:484:9  */
  assign n23697_o = n23599_o ? n23665_o : n23676_o;
  /* mmu.vhdl:481:9  */
  assign n23698_o = n23594_o ? n23696_o : n23697_o;
  /* mmu.vhdl:478:9  */
  assign n23700_o = n23580_o ? n23686_o : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* mmu.vhdl:478:9  */
  assign n23701_o = n23580_o ? n23691_o : n23698_o;
  /* mmu.vhdl:475:9  */
  assign n23703_o = n23589_o ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n23700_o;
  /* mmu.vhdl:475:9  */
  assign n23704_o = n23589_o ? n23688_o : n23701_o;
  /* mmu.vhdl:492:25  */
  assign n23705_o = r[169];
  /* mmu.vhdl:493:24  */
  assign n23706_o = r[170];
  /* mmu.vhdl:494:28  */
  assign n23707_o = r[497];
  /* mmu.vhdl:495:28  */
  assign n23708_o = r[498];
  /* mmu.vhdl:496:27  */
  assign n23709_o = r[499];
  /* mmu.vhdl:497:31  */
  assign n23710_o = r[500];
  /* mmu.vhdl:498:29  */
  assign n23711_o = r[501];
  /* mmu.vhdl:502:26  */
  assign n23712_o = r[68];
  /* mmu.vhdl:509:26  */
  assign n23713_o = r[68];
  /* mmu.vhdl:89:9  */
  always @(posedge clk)
    n23721_q <= n22495_o;
  /* mmu.vhdl:89:9  */
  assign n23722_o = {n22447_o, n23711_o, n23710_o, n23709_o, n23708_o, n23707_o, n23706_o, n23705_o};
  assign n23723_o = {n23703_o, n23704_o, n23580_o, n23712_o, n23589_o, n23575_o};
  assign n23724_o = {n23703_o, n23704_o, n23713_o, n23589_o, n23584_o};
endmodule

module loadstore1_0_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clk,
   input  rst,
   input  l_in_valid,
   input  [5:0] l_in_op,
   input  [63:0] l_in_nia,
   input  [31:0] l_in_insn,
   input  [2:0] l_in_instr_tag,
   input  [63:0] l_in_addr1,
   input  [63:0] l_in_addr2,
   input  [63:0] l_in_data,
   input  [6:0] l_in_write_reg,
   input  [3:0] l_in_length,
   input  l_in_ci,
   input  l_in_byte_reverse,
   input  l_in_sign_extend,
   input  l_in_update,
   input  [4:0] l_in_xerc,
   input  l_in_reserve,
   input  l_in_rc,
   input  l_in_virt_mode,
   input  l_in_priv_mode,
   input  l_in_mode_32bit,
   input  l_in_is_32bit,
   input  l_in_repeat,
   input  l_in_second,
   input  [63:0] l_in_msr,
   input  d_in_valid,
   input  [63:0] d_in_data,
   input  d_in_store_done,
   input  d_in_error,
   input  d_in_cache_paradox,
   input  m_in_done,
   input  m_in_err,
   input  m_in_invalid,
   input  m_in_badtree,
   input  m_in_segerr,
   input  m_in_perm_error,
   input  m_in_rc_error,
   input  [63:0] m_in_sprval,
   input  dc_stall,
   output e_out_busy,
   output e_out_in_progress,
   output e_out_interrupt,
   output l_out_valid,
   output [2:0] l_out_instr_tag,
   output l_out_write_enable,
   output [6:0] l_out_write_reg,
   output [63:0] l_out_write_data,
   output [4:0] l_out_xerc,
   output l_out_rc,
   output l_out_store_done,
   output l_out_interrupt,
   output [11:0] l_out_intr_vec,
   output [63:0] l_out_srr0,
   output [15:0] l_out_srr1,
   output d_out_valid,
   output d_out_hold,
   output d_out_load,
   output d_out_dcbz,
   output d_out_nc,
   output d_out_reserve,
   output d_out_atomic,
   output d_out_atomic_last,
   output d_out_virt_mode,
   output d_out_priv_mode,
   output [63:0] d_out_addr,
   output [63:0] d_out_data,
   output [7:0] d_out_byte_sel,
   output m_out_valid,
   output m_out_tlbie,
   output m_out_slbia,
   output m_out_mtspr,
   output m_out_iside,
   output m_out_load,
   output m_out_priv,
   output [9:0] m_out_sprn,
   output [63:0] m_out_addr,
   output [63:0] m_out_rs,
   output events_load_complete,
   output events_store_complete,
   output events_itlb_miss,
   output [9:0] log_out);
  wire [389:0] n19326_o;
  wire n19328_o;
  wire n19329_o;
  wire n19330_o;
  wire n19332_o;
  wire [2:0] n19333_o;
  wire n19334_o;
  wire [6:0] n19335_o;
  wire [63:0] n19336_o;
  wire [4:0] n19337_o;
  wire n19338_o;
  wire n19339_o;
  wire n19340_o;
  wire [11:0] n19341_o;
  wire [63:0] n19342_o;
  wire [15:0] n19343_o;
  wire n19345_o;
  wire n19346_o;
  wire n19347_o;
  wire n19348_o;
  wire n19349_o;
  wire n19350_o;
  wire n19351_o;
  wire n19352_o;
  wire n19353_o;
  wire n19354_o;
  wire [63:0] n19355_o;
  wire [63:0] n19356_o;
  wire [7:0] n19357_o;
  wire [67:0] n19358_o;
  wire n19360_o;
  wire n19361_o;
  wire n19362_o;
  wire n19363_o;
  wire n19364_o;
  wire n19365_o;
  wire n19366_o;
  wire [9:0] n19367_o;
  wire [63:0] n19368_o;
  wire [63:0] n19369_o;
  wire [70:0] n19370_o;
  wire n19372_o;
  wire n19373_o;
  wire n19374_o;
  wire [272:0] req_in;
  wire [337:0] r1;
  wire [337:0] r1in;
  wire [373:0] r2;
  wire [373:0] r2in;
  wire [380:0] r3;
  wire [380:0] r3in;
  wire busy;
  wire complete;
  wire in_progress;
  wire flushing;
  wire [31:0] store_sp_data;
  wire [63:0] load_dp_data;
  wire [63:0] store_data;
  wire stage1_issue_enable;
  wire [272:0] stage1_req;
  wire stage1_dcreq;
  wire stage1_dreq;
  wire stage2_busy_next;
  wire stage3_busy_next;
  wire [272:0] n19390_o;
  wire n19391_o;
  wire [272:0] n19392_o;
  wire n19393_o;
  wire n19394_o;
  wire n19395_o;
  wire n19396_o;
  wire n19397_o;
  wire n19398_o;
  wire n19399_o;
  wire n19400_o;
  wire [336:0] n19401_o;
  wire [336:0] n19402_o;
  wire [336:0] n19403_o;
  wire [2:0] n19404_o;
  wire n19405_o;
  wire n19406_o;
  wire [303:0] n19407_o;
  wire [303:0] n19408_o;
  wire [303:0] n19409_o;
  wire [2:0] n19410_o;
  wire [2:0] n19411_o;
  wire [65:0] n19412_o;
  wire [65:0] n19413_o;
  wire [65:0] n19414_o;
  wire [95:0] n19415_o;
  wire [1:0] n19416_o;
  wire [1:0] n19417_o;
  wire [1:0] n19418_o;
  wire [2:0] n19419_o;
  wire [2:0] n19420_o;
  wire [2:0] n19421_o;
  wire n19422_o;
  wire n19423_o;
  wire [77:0] n19424_o;
  wire [77:0] n19425_o;
  wire [77:0] n19426_o;
  wire n19427_o;
  wire n19428_o;
  wire [63:0] n19429_o;
  wire [63:0] n19430_o;
  wire [63:0] n19431_o;
  wire [95:0] n19432_o;
  wire [95:0] n19433_o;
  wire [38:0] n19434_o;
  wire [38:0] n19435_o;
  wire [38:0] n19436_o;
  wire [1:0] n19437_o;
  wire [1:0] n19438_o;
  wire [94:0] n19439_o;
  wire [94:0] n19440_o;
  wire [94:0] n19441_o;
  wire n19443_o;
  wire [337:0] n19449_o;
  wire [373:0] n19451_o;
  wire [380:0] n19453_o;
  wire n19462_o;
  localparam [30:0] n19463_o = 31'b0000000000000000000000000000000;
  wire [10:0] n19464_o;
  wire n19466_o;
  wire n19467_o;
  wire [29:0] n19468_o;
  wire n19470_o;
  wire [21:0] n19471_o;
  wire [22:0] n19473_o;
  wire [4:0] n19474_o;
  wire [4:0] n19476_o;
  wire [1:0] n19484_o;
  wire n19486_o;
  wire [21:0] n19487_o;
  wire [22:0] n19489_o;
  wire n19491_o;
  wire [20:0] n19492_o;
  wire [22:0] n19494_o;
  wire n19496_o;
  wire [19:0] n19497_o;
  wire [22:0] n19499_o;
  wire [2:0] n19500_o;
  reg [22:0] n19501_o;
  wire [2:0] n19503_o;
  wire n19505_o;
  wire [18:0] n19506_o;
  wire [22:0] n19508_o;
  wire n19510_o;
  wire [14:0] n19511_o;
  wire [22:0] n19513_o;
  wire n19515_o;
  wire [10:0] n19516_o;
  wire [22:0] n19518_o;
  wire n19520_o;
  wire [6:0] n19521_o;
  wire [22:0] n19523_o;
  wire n19525_o;
  wire [2:0] n19526_o;
  wire [22:0] n19528_o;
  wire [4:0] n19529_o;
  reg [22:0] n19530_o;
  wire [22:0] n19532_o;
  wire [22:0] n19533_o;
  wire [30:0] n19536_o;
  wire [22:0] n19537_o;
  wire [22:0] n19538_o;
  wire [7:0] n19539_o;
  wire [7:0] n19540_o;
  wire [7:0] n19541_o;
  wire [22:0] n19555_o;
  wire [7:0] n19556_o;
  wire [7:0] n19557_o;
  wire n19558_o;
  wire [7:0] n19559_o;
  wire n19560_o;
  wire [10:0] n19561_o;
  wire [10:0] n19563_o;
  wire n19564_o;
  wire n19565_o;
  wire [5:0] n19566_o;
  wire [10:0] n19567_o;
  wire [10:0] n19569_o;
  wire [4:0] n19570_o;
  wire [4:0] n19572_o;
  wire [10:0] n19574_o;
  wire [4:0] n19576_o;
  wire [10:0] n19577_o;
  wire [4:0] n19579_o;
  wire [10:0] n19581_o;
  wire [4:0] n19583_o;
  wire n19585_o;
  wire [1:0] n19593_o;
  wire n19595_o;
  wire [21:0] n19596_o;
  wire [22:0] n19598_o;
  wire n19600_o;
  wire [20:0] n19601_o;
  wire [22:0] n19603_o;
  wire n19605_o;
  wire [19:0] n19606_o;
  wire [22:0] n19608_o;
  wire [2:0] n19609_o;
  reg [22:0] n19610_o;
  wire [2:0] n19612_o;
  wire n19614_o;
  wire [18:0] n19615_o;
  wire [22:0] n19617_o;
  wire n19619_o;
  wire [14:0] n19620_o;
  wire [22:0] n19622_o;
  wire n19624_o;
  wire [10:0] n19625_o;
  wire [22:0] n19627_o;
  wire n19629_o;
  wire [6:0] n19630_o;
  wire [22:0] n19632_o;
  wire n19634_o;
  wire [2:0] n19635_o;
  wire [22:0] n19637_o;
  wire [4:0] n19638_o;
  reg [22:0] n19639_o;
  wire [31:0] n19654_o;
  wire [4:0] n19659_o;
  wire [4:0] n19660_o;
  wire [9:0] n19661_o;
  wire n19664_o;
  localparam [272:0] n19665_o = 273'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [2:0] n19667_o;
  wire n19670_o;
  wire [11:0] n19672_o;
  wire [6:0] n19673_o;
  wire [3:0] n19675_o;
  wire [3:0] n19677_o;
  wire n19679_o;
  wire n19681_o;
  wire [2:0] n19683_o;
  wire n19684_o;
  wire [4:0] n19686_o;
  wire n19688_o;
  wire n19690_o;
  wire [1:0] n19692_o;
  wire n19693_o;
  wire n19695_o;
  wire n19697_o;
  wire n19700_o;
  wire [63:0] n19701_o;
  wire [3:0] n19702_o;
  wire [63:0] n19703_o;
  wire [63:0] n19704_o;
  wire [63:0] n19705_o;
  wire n19706_o;
  wire n19708_o;
  wire [63:0] n19710_o;
  wire [63:0] n19711_o;
  wire [63:0] n19712_o;
  wire n19714_o;
  wire n19715_o;
  wire n19716_o;
  wire [60:0] n19717_o;
  wire [60:0] n19719_o;
  wire [2:0] n19720_o;
  wire [63:0] n19721_o;
  wire n19725_o;
  wire [31:0] n19727_o;
  wire [31:0] n19728_o;
  wire [31:0] n19729_o;
  wire [31:0] n19730_o;
  wire [31:0] n19731_o;
  wire [31:0] n19732_o;
  wire [31:0] n19733_o;
  wire [31:0] n19734_o;
  wire [31:0] n19735_o;
  wire [31:0] n19736_o;
  wire [31:0] n19737_o;
  wire [63:0] n19738_o;
  wire [15:0] n19739_o;
  wire [63:0] n19740_o;
  wire [3:0] n19741_o;
  wire n19743_o;
  wire n19744_o;
  wire n19745_o;
  wire n19746_o;
  wire n19748_o;
  wire [2:0] n19749_o;
  wire [2:0] n19751_o;
  wire [272:0] n19753_o;
  wire [3:0] n19754_o;
  wire [63:0] n19755_o;
  wire [2:0] n19756_o;
  wire n19769_o;
  wire n19772_o;
  wire n19775_o;
  wire n19778_o;
  wire [3:0] n19780_o;
  reg [7:0] n19781_o;
  wire [15:0] n19783_o;
  wire [30:0] n19785_o;
  wire [15:0] n19786_o;
  wire [7:0] n19787_o;
  wire [7:0] n19789_o;
  wire [7:0] n19790_o;
  wire n19792_o;
  wire n19794_o;
  wire n19795_o;
  wire [63:0] n19797_o;
  wire [2:0] n19798_o;
  wire [2:0] n19799_o;
  wire n19800_o;
  wire n19801_o;
  wire n19802_o;
  wire n19803_o;
  wire n19804_o;
  wire n19805_o;
  wire n19806_o;
  wire n19807_o;
  wire n19808_o;
  wire n19809_o;
  wire n19810_o;
  wire n19811_o;
  wire [63:0] n19812_o;
  wire n19813_o;
  wire n19814_o;
  wire n19815_o;
  wire [5:0] n19816_o;
  wire n19818_o;
  wire n19819_o;
  wire n19820_o;
  wire n19821_o;
  wire n19822_o;
  wire n19824_o;
  wire n19825_o;
  wire n19827_o;
  wire n19828_o;
  wire n19830_o;
  wire n19831_o;
  wire n19832_o;
  wire n19833_o;
  wire n19834_o;
  wire n19835_o;
  wire [5:0] n19836_o;
  wire n19839_o;
  wire n19840_o;
  wire n19841_o;
  wire n19842_o;
  wire n19843_o;
  wire n19844_o;
  wire n19846_o;
  wire n19848_o;
  wire n19850_o;
  wire n19852_o;
  wire n19853_o;
  wire n19854_o;
  wire n19855_o;
  wire n19856_o;
  wire n19858_o;
  wire [3:0] n19860_o;
  wire [6:0] n19861_o;
  wire [272:0] n19862_o;
  wire n19863_o;
  wire n19865_o;
  wire [63:0] n19867_o;
  wire n19868_o;
  wire n19871_o;
  wire n19874_o;
  wire n19876_o;
  wire n19877_o;
  wire n19878_o;
  wire n19880_o;
  wire [63:0] n19882_o;
  wire n19885_o;
  wire [6:0] n19886_o;
  wire n19887_o;
  reg n19888_o;
  wire n19889_o;
  reg n19890_o;
  wire n19891_o;
  reg n19892_o;
  wire n19893_o;
  reg n19894_o;
  wire n19895_o;
  reg n19896_o;
  wire n19897_o;
  reg n19898_o;
  wire n19899_o;
  reg n19900_o;
  wire n19901_o;
  reg n19902_o;
  wire n19903_o;
  reg n19904_o;
  reg [63:0] n19905_o;
  reg n19906_o;
  reg n19907_o;
  reg n19908_o;
  wire n19910_o;
  wire n19918_o;
  wire n19919_o;
  wire n19920_o;
  wire [272:0] n19921_o;
  wire n19922_o;
  wire [272:0] n19923_o;
  wire n19924_o;
  wire n19925_o;
  wire [272:0] n19926_o;
  wire n19927_o;
  wire n19928_o;
  wire n19929_o;
  wire [272:0] n19930_o;
  wire n19931_o;
  wire n19932_o;
  wire n19933_o;
  wire [272:0] n19934_o;
  wire n19935_o;
  wire [272:0] n19936_o;
  wire [2:0] n19937_o;
  wire [2:0] n19939_o;
  wire [2:0] n19941_o;
  wire [272:0] n19943_o;
  wire [272:0] n19948_o;
  wire n19949_o;
  wire [272:0] n19950_o;
  wire n19951_o;
  wire n19952_o;
  wire n19953_o;
  wire n19954_o;
  wire n19955_o;
  wire n19956_o;
  wire n19957_o;
  wire n19958_o;
  wire n19959_o;
  wire [272:0] n19960_o;
  wire n19961_o;
  wire [272:0] n19962_o;
  wire n19963_o;
  wire n19964_o;
  wire [272:0] n19965_o;
  wire n19966_o;
  wire n19967_o;
  wire n19968_o;
  wire n19969_o;
  wire n19970_o;
  wire n19971_o;
  wire n19972_o;
  wire n19973_o;
  wire n19974_o;
  wire n19975_o;
  wire n19976_o;
  wire n19977_o;
  wire n19978_o;
  wire n19979_o;
  wire n19980_o;
  wire n19981_o;
  wire [272:0] n19982_o;
  wire n19983_o;
  wire [272:0] n19984_o;
  wire n19985_o;
  wire n19986_o;
  wire n19987_o;
  wire n19988_o;
  wire n19989_o;
  wire [272:0] n19990_o;
  wire n19991_o;
  wire [272:0] n19992_o;
  wire n19993_o;
  wire n19994_o;
  wire n19995_o;
  wire n19996_o;
  wire [272:0] n19997_o;
  wire n19998_o;
  wire [272:0] n19999_o;
  wire n20000_o;
  wire n20001_o;
  wire n20002_o;
  wire n20003_o;
  wire n20009_o;
  wire n20012_o;
  wire n20013_o;
  wire [270:0] n20014_o;
  wire n20015_o;
  wire n20016_o;
  wire [272:0] n20017_o;
  wire n20018_o;
  wire n20019_o;
  wire n20020_o;
  wire [272:0] n20021_o;
  wire [63:0] n20022_o;
  wire [63:0] n20023_o;
  wire [63:0] n20024_o;
  wire [64:0] n20026_o;
  wire [272:0] n20030_o;
  wire n20033_o;
  wire [272:0] n20035_o;
  wire n20036_o;
  wire [272:0] n20037_o;
  wire n20038_o;
  wire n20039_o;
  wire n20040_o;
  wire n20041_o;
  wire n20042_o;
  wire n20043_o;
  wire n20044_o;
  wire n20046_o;
  wire [272:0] n20047_o;
  wire n20048_o;
  wire [272:0] n20049_o;
  wire n20050_o;
  wire n20051_o;
  wire [272:0] n20052_o;
  wire n20053_o;
  wire n20054_o;
  wire n20055_o;
  wire [60:0] n20057_o;
  wire [60:0] n20059_o;
  wire [63:0] n20061_o;
  wire [272:0] n20062_o;
  wire n20063_o;
  wire n20065_o;
  wire n20066_o;
  wire [30:0] n20067_o;
  wire [31:0] n20068_o;
  wire [272:0] n20069_o;
  wire [7:0] n20070_o;
  wire [71:0] n20071_o;
  wire [71:0] n20072_o;
  wire [71:0] n20073_o;
  wire [71:0] n20074_o;
  wire [71:0] n20075_o;
  wire n20076_o;
  wire n20077_o;
  wire n20078_o;
  wire n20079_o;
  wire n20081_o;
  wire [71:0] n20082_o;
  wire [71:0] n20083_o;
  wire [71:0] n20084_o;
  wire [71:0] n20085_o;
  wire n20086_o;
  wire n20087_o;
  wire n20088_o;
  wire n20089_o;
  wire n20090_o;
  wire n20091_o;
  wire n20092_o;
  wire n20093_o;
  wire n20094_o;
  wire [71:0] n20095_o;
  wire [71:0] n20096_o;
  wire [71:0] n20097_o;
  wire [71:0] n20098_o;
  wire n20099_o;
  wire n20100_o;
  wire n20101_o;
  wire n20102_o;
  wire n20103_o;
  wire n20104_o;
  wire n20105_o;
  wire n20106_o;
  wire n20107_o;
  wire [71:0] n20108_o;
  wire [71:0] n20109_o;
  wire [71:0] n20110_o;
  wire [71:0] n20111_o;
  wire n20112_o;
  wire n20113_o;
  wire n20114_o;
  wire n20115_o;
  wire n20117_o;
  wire n20118_o;
  wire n20119_o;
  wire n20120_o;
  wire n20121_o;
  wire [63:0] n20122_o;
  wire [63:0] n20123_o;
  wire [63:0] n20124_o;
  wire [71:0] n20125_o;
  wire [71:0] n20126_o;
  wire [71:0] n20127_o;
  wire [71:0] n20128_o;
  wire n20129_o;
  wire n20130_o;
  wire n20131_o;
  wire n20132_o;
  wire [64:0] n20139_o;
  wire [64:0] n20140_o;
  wire [64:0] n20141_o;
  wire [120:0] n20142_o;
  wire [120:0] n20143_o;
  wire [120:0] n20144_o;
  wire n20145_o;
  wire n20146_o;
  wire n20148_o;
  wire n20149_o;
  wire n20150_o;
  wire n20151_o;
  wire [12:0] n20152_o;
  wire [12:0] n20153_o;
  wire [12:0] n20154_o;
  wire n20156_o;
  wire [272:0] n20157_o;
  wire n20158_o;
  wire n20159_o;
  wire n20160_o;
  wire n20161_o;
  wire n20162_o;
  wire n20163_o;
  wire n20164_o;
  wire [272:0] n20165_o;
  wire [337:0] n20166_o;
  wire [2:0] n20177_o;
  wire [2:0] n20179_o;
  wire [272:0] n20180_o;
  wire [2:0] n20181_o;
  wire [2:0] n20182_o;
  wire [2:0] n20192_o;
  wire [272:0] n20193_o;
  wire [2:0] n20194_o;
  wire [2:0] n20195_o;
  wire [2:0] n20205_o;
  wire [272:0] n20206_o;
  wire [2:0] n20207_o;
  wire [2:0] n20208_o;
  wire [2:0] n20218_o;
  wire [272:0] n20219_o;
  wire [2:0] n20220_o;
  wire [2:0] n20221_o;
  wire [2:0] n20231_o;
  wire [272:0] n20232_o;
  wire [2:0] n20233_o;
  wire [2:0] n20234_o;
  wire [2:0] n20244_o;
  wire [272:0] n20245_o;
  wire [2:0] n20246_o;
  wire [2:0] n20247_o;
  wire [2:0] n20257_o;
  wire [272:0] n20258_o;
  wire [2:0] n20259_o;
  wire [2:0] n20260_o;
  wire [2:0] n20270_o;
  wire [272:0] n20271_o;
  wire [2:0] n20272_o;
  wire [2:0] n20273_o;
  wire n20282_o;
  wire [272:0] n20283_o;
  wire n20284_o;
  wire n20285_o;
  wire n20286_o;
  wire n20287_o;
  wire [272:0] n20288_o;
  wire n20289_o;
  wire n20290_o;
  wire n20291_o;
  wire n20292_o;
  wire [63:0] n20294_o;
  wire [114:0] n20295_o;
  wire [93:0] n20296_o;
  wire [272:0] n20297_o;
  wire n20298_o;
  wire [272:0] n20299_o;
  wire n20300_o;
  wire n20301_o;
  wire [272:0] n20302_o;
  wire n20303_o;
  wire n20304_o;
  wire n20305_o;
  wire [272:0] n20306_o;
  wire n20307_o;
  wire [272:0] n20308_o;
  wire n20309_o;
  wire n20310_o;
  wire n20311_o;
  wire n20312_o;
  wire n20313_o;
  wire [272:0] n20314_o;
  wire n20315_o;
  wire [272:0] n20316_o;
  wire n20317_o;
  wire n20318_o;
  wire [272:0] n20319_o;
  wire n20320_o;
  wire [272:0] n20321_o;
  wire n20322_o;
  wire [272:0] n20323_o;
  wire n20324_o;
  wire n20325_o;
  wire [272:0] n20326_o;
  wire n20327_o;
  wire [272:0] n20328_o;
  wire n20329_o;
  wire n20330_o;
  wire n20331_o;
  wire n20332_o;
  wire [272:0] n20333_o;
  wire n20334_o;
  wire n20335_o;
  wire [272:0] n20336_o;
  wire n20337_o;
  wire n20338_o;
  wire n20339_o;
  wire [272:0] n20340_o;
  wire n20341_o;
  wire [272:0] n20343_o;
  wire n20344_o;
  wire [272:0] n20345_o;
  wire n20346_o;
  wire n20347_o;
  wire [272:0] n20349_o;
  wire n20350_o;
  wire [1:0] n20353_o;
  wire [1:0] n20354_o;
  wire [1:0] n20355_o;
  wire [272:0] n20356_o;
  wire [2:0] n20357_o;
  wire [2:0] n20359_o;
  wire [3:0] n20361_o;
  wire [3:0] n20363_o;
  wire [3:0] n20364_o;
  wire n20365_o;
  wire [2:0] n20366_o;
  wire [272:0] n20367_o;
  wire [2:0] n20368_o;
  wire [2:0] n20370_o;
  wire [3:0] n20372_o;
  wire [3:0] n20374_o;
  wire [3:0] n20375_o;
  wire n20376_o;
  wire [2:0] n20377_o;
  wire [272:0] n20378_o;
  wire [2:0] n20379_o;
  wire [2:0] n20381_o;
  wire [3:0] n20383_o;
  wire [3:0] n20385_o;
  wire [3:0] n20386_o;
  wire n20387_o;
  wire [2:0] n20388_o;
  wire [272:0] n20389_o;
  wire [2:0] n20390_o;
  wire [2:0] n20392_o;
  wire [3:0] n20394_o;
  wire [3:0] n20396_o;
  wire [3:0] n20397_o;
  wire n20398_o;
  wire [2:0] n20399_o;
  wire [272:0] n20400_o;
  wire [2:0] n20401_o;
  wire [2:0] n20403_o;
  wire [3:0] n20405_o;
  wire [3:0] n20407_o;
  wire [3:0] n20408_o;
  wire n20409_o;
  wire [2:0] n20410_o;
  wire [272:0] n20411_o;
  wire [2:0] n20412_o;
  wire [2:0] n20414_o;
  wire [3:0] n20416_o;
  wire [3:0] n20418_o;
  wire [3:0] n20419_o;
  wire n20420_o;
  wire [2:0] n20421_o;
  wire [272:0] n20422_o;
  wire [2:0] n20423_o;
  wire [2:0] n20425_o;
  wire [3:0] n20427_o;
  wire [3:0] n20429_o;
  wire [3:0] n20430_o;
  wire n20431_o;
  wire [2:0] n20432_o;
  wire [272:0] n20433_o;
  wire [2:0] n20434_o;
  wire [2:0] n20436_o;
  wire [3:0] n20438_o;
  wire [3:0] n20440_o;
  wire [3:0] n20441_o;
  wire n20442_o;
  wire [2:0] n20443_o;
  wire n20444_o;
  wire [1:0] n20448_o;
  wire n20449_o;
  wire n20450_o;
  wire [1:0] n20451_o;
  wire [1:0] n20452_o;
  wire [373:0] n20453_o;
  wire n20454_o;
  wire n20455_o;
  wire [303:0] n20456_o;
  wire [303:0] n20457_o;
  wire [303:0] n20458_o;
  wire [1:0] n20459_o;
  wire [1:0] n20460_o;
  wire [66:0] n20461_o;
  wire [66:0] n20462_o;
  wire [66:0] n20463_o;
  wire [272:0] n20469_o;
  wire n20470_o;
  wire n20471_o;
  wire n20472_o;
  wire n20474_o;
  wire [373:0] n20475_o;
  localparam [15:0] n20500_o = 16'b0000000000000000;
  localparam [2:0] n20503_o = 3'b000;
  wire [2:0] n20504_o;
  wire [2:0] n20513_o;
  wire [2:0] n20522_o;
  wire [2:0] n20531_o;
  wire [2:0] n20540_o;
  wire [2:0] n20549_o;
  wire [2:0] n20558_o;
  wire [2:0] n20567_o;
  wire [272:0] n20576_o;
  wire n20577_o;
  wire [272:0] n20578_o;
  wire n20579_o;
  wire n20580_o;
  wire n20581_o;
  wire n20582_o;
  wire n20583_o;
  wire n20584_o;
  wire n20585_o;
  wire n20586_o;
  wire n20587_o;
  wire n20588_o;
  wire n20589_o;
  wire n20590_o;
  wire n20591_o;
  wire n20592_o;
  wire n20593_o;
  wire n20594_o;
  wire n20595_o;
  wire n20596_o;
  wire [63:0] n20597_o;
  wire n20598_o;
  wire n20599_o;
  wire n20600_o;
  wire [63:0] n20601_o;
  wire n20602_o;
  wire n20603_o;
  wire n20604_o;
  wire n20605_o;
  wire [63:0] n20606_o;
  wire n20607_o;
  wire n20608_o;
  wire n20609_o;
  wire n20610_o;
  wire [63:0] n20611_o;
  wire n20612_o;
  wire n20613_o;
  wire n20614_o;
  wire n20615_o;
  wire [272:0] n20616_o;
  wire [3:0] n20617_o;
  wire [30:0] n20618_o;
  wire [31:0] n20619_o;
  wire n20621_o;
  wire [272:0] n20622_o;
  wire n20623_o;
  wire n20624_o;
  wire n20625_o;
  wire [1:0] n20627_o;
  wire [1:0] n20629_o;
  wire [1:0] n20631_o;
  wire [272:0] n20632_o;
  wire [3:0] n20633_o;
  wire [30:0] n20634_o;
  wire [31:0] n20635_o;
  wire n20637_o;
  wire [272:0] n20638_o;
  wire n20639_o;
  wire n20640_o;
  wire n20641_o;
  wire [1:0] n20643_o;
  wire [1:0] n20645_o;
  wire [1:0] n20647_o;
  wire [272:0] n20648_o;
  wire [3:0] n20649_o;
  wire [30:0] n20650_o;
  wire [31:0] n20651_o;
  wire n20653_o;
  wire [272:0] n20654_o;
  wire n20655_o;
  wire n20656_o;
  wire n20657_o;
  wire [1:0] n20659_o;
  wire [1:0] n20661_o;
  wire [1:0] n20663_o;
  wire [272:0] n20664_o;
  wire [3:0] n20665_o;
  wire [30:0] n20666_o;
  wire [31:0] n20667_o;
  wire n20669_o;
  wire [272:0] n20670_o;
  wire n20671_o;
  wire n20672_o;
  wire n20673_o;
  wire [1:0] n20675_o;
  wire [1:0] n20677_o;
  wire [1:0] n20679_o;
  wire [272:0] n20680_o;
  wire [3:0] n20681_o;
  wire [30:0] n20682_o;
  wire [31:0] n20683_o;
  wire n20685_o;
  wire [272:0] n20686_o;
  wire n20687_o;
  wire n20688_o;
  wire n20689_o;
  wire [1:0] n20691_o;
  wire [1:0] n20693_o;
  wire [1:0] n20695_o;
  wire [272:0] n20696_o;
  wire [3:0] n20697_o;
  wire [30:0] n20698_o;
  wire [31:0] n20699_o;
  wire n20701_o;
  wire [272:0] n20702_o;
  wire n20703_o;
  wire n20704_o;
  wire n20705_o;
  wire [1:0] n20707_o;
  wire [1:0] n20709_o;
  wire [1:0] n20711_o;
  wire [272:0] n20712_o;
  wire [3:0] n20713_o;
  wire [30:0] n20714_o;
  wire [31:0] n20715_o;
  wire n20717_o;
  wire [272:0] n20718_o;
  wire n20719_o;
  wire n20720_o;
  wire n20721_o;
  wire [1:0] n20723_o;
  wire [1:0] n20725_o;
  wire [1:0] n20727_o;
  wire [272:0] n20728_o;
  wire [3:0] n20729_o;
  wire [30:0] n20730_o;
  wire [31:0] n20731_o;
  wire n20733_o;
  wire [272:0] n20734_o;
  wire n20735_o;
  wire n20736_o;
  wire n20737_o;
  wire [1:0] n20739_o;
  wire [1:0] n20741_o;
  wire [1:0] n20743_o;
  wire [15:0] n20744_o;
  wire [1:0] n20745_o;
  wire [7:0] n20746_o;
  wire n20748_o;
  wire [63:0] n20749_o;
  wire [7:0] n20750_o;
  wire n20752_o;
  wire [272:0] n20753_o;
  wire n20754_o;
  wire n20755_o;
  wire [272:0] n20756_o;
  wire n20757_o;
  wire n20758_o;
  wire [272:0] n20759_o;
  wire n20760_o;
  wire n20761_o;
  wire [272:0] n20762_o;
  wire n20763_o;
  wire n20764_o;
  wire [272:0] n20765_o;
  wire n20766_o;
  wire n20767_o;
  wire [272:0] n20768_o;
  wire n20769_o;
  wire n20770_o;
  wire [272:0] n20771_o;
  wire n20772_o;
  wire n20773_o;
  wire [272:0] n20774_o;
  wire n20775_o;
  wire n20776_o;
  wire [3:0] n20777_o;
  wire [3:0] n20778_o;
  wire [7:0] n20779_o;
  wire [1:0] n20780_o;
  reg [7:0] n20781_o;
  wire [15:0] n20782_o;
  wire [1:0] n20783_o;
  wire [7:0] n20784_o;
  wire n20786_o;
  wire [63:0] n20787_o;
  wire [7:0] n20788_o;
  wire n20790_o;
  wire [272:0] n20791_o;
  wire n20792_o;
  wire n20793_o;
  wire [272:0] n20794_o;
  wire n20795_o;
  wire n20796_o;
  wire [272:0] n20797_o;
  wire n20798_o;
  wire n20799_o;
  wire [272:0] n20800_o;
  wire n20801_o;
  wire n20802_o;
  wire [272:0] n20803_o;
  wire n20804_o;
  wire n20805_o;
  wire [272:0] n20806_o;
  wire n20807_o;
  wire n20808_o;
  wire [272:0] n20809_o;
  wire n20810_o;
  wire n20811_o;
  wire [272:0] n20812_o;
  wire n20813_o;
  wire n20814_o;
  wire [3:0] n20815_o;
  wire [3:0] n20816_o;
  wire [7:0] n20817_o;
  wire [1:0] n20818_o;
  reg [7:0] n20819_o;
  wire [15:0] n20820_o;
  wire [1:0] n20821_o;
  wire [7:0] n20822_o;
  wire n20824_o;
  wire [63:0] n20825_o;
  wire [7:0] n20826_o;
  wire n20828_o;
  wire [272:0] n20829_o;
  wire n20830_o;
  wire n20831_o;
  wire [272:0] n20832_o;
  wire n20833_o;
  wire n20834_o;
  wire [272:0] n20835_o;
  wire n20836_o;
  wire n20837_o;
  wire [272:0] n20838_o;
  wire n20839_o;
  wire n20840_o;
  wire [272:0] n20841_o;
  wire n20842_o;
  wire n20843_o;
  wire [272:0] n20844_o;
  wire n20845_o;
  wire n20846_o;
  wire [272:0] n20847_o;
  wire n20848_o;
  wire n20849_o;
  wire [272:0] n20850_o;
  wire n20851_o;
  wire n20852_o;
  wire [3:0] n20853_o;
  wire [3:0] n20854_o;
  wire [7:0] n20855_o;
  wire [1:0] n20856_o;
  reg [7:0] n20857_o;
  wire [15:0] n20858_o;
  wire [1:0] n20859_o;
  wire [7:0] n20860_o;
  wire n20862_o;
  wire [63:0] n20863_o;
  wire [7:0] n20864_o;
  wire n20866_o;
  wire [272:0] n20867_o;
  wire n20868_o;
  wire n20869_o;
  wire [272:0] n20870_o;
  wire n20871_o;
  wire n20872_o;
  wire [272:0] n20873_o;
  wire n20874_o;
  wire n20875_o;
  wire [272:0] n20876_o;
  wire n20877_o;
  wire n20878_o;
  wire [272:0] n20879_o;
  wire n20880_o;
  wire n20881_o;
  wire [272:0] n20882_o;
  wire n20883_o;
  wire n20884_o;
  wire [272:0] n20885_o;
  wire n20886_o;
  wire n20887_o;
  wire [272:0] n20888_o;
  wire n20889_o;
  wire n20890_o;
  wire [3:0] n20891_o;
  wire [3:0] n20892_o;
  wire [7:0] n20893_o;
  wire [1:0] n20894_o;
  reg [7:0] n20895_o;
  wire [15:0] n20896_o;
  wire [1:0] n20897_o;
  wire [7:0] n20898_o;
  wire n20900_o;
  wire [63:0] n20901_o;
  wire [7:0] n20902_o;
  wire n20904_o;
  wire [272:0] n20905_o;
  wire n20906_o;
  wire n20907_o;
  wire [272:0] n20908_o;
  wire n20909_o;
  wire n20910_o;
  wire [272:0] n20911_o;
  wire n20912_o;
  wire n20913_o;
  wire [272:0] n20914_o;
  wire n20915_o;
  wire n20916_o;
  wire [272:0] n20917_o;
  wire n20918_o;
  wire n20919_o;
  wire [272:0] n20920_o;
  wire n20921_o;
  wire n20922_o;
  wire [272:0] n20923_o;
  wire n20924_o;
  wire n20925_o;
  wire [272:0] n20926_o;
  wire n20927_o;
  wire n20928_o;
  wire [3:0] n20929_o;
  wire [3:0] n20930_o;
  wire [7:0] n20931_o;
  wire [1:0] n20932_o;
  reg [7:0] n20933_o;
  wire [15:0] n20934_o;
  wire [1:0] n20935_o;
  wire [7:0] n20936_o;
  wire n20938_o;
  wire [63:0] n20939_o;
  wire [7:0] n20940_o;
  wire n20942_o;
  wire [272:0] n20943_o;
  wire n20944_o;
  wire n20945_o;
  wire [272:0] n20946_o;
  wire n20947_o;
  wire n20948_o;
  wire [272:0] n20949_o;
  wire n20950_o;
  wire n20951_o;
  wire [272:0] n20952_o;
  wire n20953_o;
  wire n20954_o;
  wire [272:0] n20955_o;
  wire n20956_o;
  wire n20957_o;
  wire [272:0] n20958_o;
  wire n20959_o;
  wire n20960_o;
  wire [272:0] n20961_o;
  wire n20962_o;
  wire n20963_o;
  wire [272:0] n20964_o;
  wire n20965_o;
  wire n20966_o;
  wire [3:0] n20967_o;
  wire [3:0] n20968_o;
  wire [7:0] n20969_o;
  wire [1:0] n20970_o;
  reg [7:0] n20971_o;
  wire [15:0] n20972_o;
  wire [1:0] n20973_o;
  wire [7:0] n20974_o;
  wire n20976_o;
  wire [63:0] n20977_o;
  wire [7:0] n20978_o;
  wire n20980_o;
  wire [272:0] n20981_o;
  wire n20982_o;
  wire n20983_o;
  wire [272:0] n20984_o;
  wire n20985_o;
  wire n20986_o;
  wire [272:0] n20987_o;
  wire n20988_o;
  wire n20989_o;
  wire [272:0] n20990_o;
  wire n20991_o;
  wire n20992_o;
  wire [272:0] n20993_o;
  wire n20994_o;
  wire n20995_o;
  wire [272:0] n20996_o;
  wire n20997_o;
  wire n20998_o;
  wire [272:0] n20999_o;
  wire n21000_o;
  wire n21001_o;
  wire [272:0] n21002_o;
  wire n21003_o;
  wire n21004_o;
  wire [3:0] n21005_o;
  wire [3:0] n21006_o;
  wire [7:0] n21007_o;
  wire [1:0] n21008_o;
  reg [7:0] n21009_o;
  wire [15:0] n21010_o;
  wire [1:0] n21011_o;
  wire [7:0] n21012_o;
  wire n21014_o;
  wire [63:0] n21015_o;
  wire [7:0] n21016_o;
  wire n21018_o;
  wire [272:0] n21019_o;
  wire n21020_o;
  wire n21021_o;
  wire [272:0] n21022_o;
  wire n21023_o;
  wire n21024_o;
  wire [272:0] n21025_o;
  wire n21026_o;
  wire n21027_o;
  wire [272:0] n21028_o;
  wire n21029_o;
  wire n21030_o;
  wire [272:0] n21031_o;
  wire n21032_o;
  wire n21033_o;
  wire [272:0] n21034_o;
  wire n21035_o;
  wire n21036_o;
  wire [272:0] n21037_o;
  wire n21038_o;
  wire n21039_o;
  wire [272:0] n21040_o;
  wire n21041_o;
  wire n21042_o;
  wire [3:0] n21043_o;
  wire [3:0] n21044_o;
  wire [7:0] n21045_o;
  wire [1:0] n21046_o;
  reg [7:0] n21047_o;
  wire [63:0] n21048_o;
  wire [31:0] n21049_o;
  wire [63:0] n21052_o;
  wire [22:0] n21053_o;
  wire n21054_o;
  wire [63:0] n21057_o;
  wire [22:0] n21058_o;
  wire n21070_o;
  wire n21073_o;
  wire n21075_o;
  wire n21077_o;
  wire n21079_o;
  wire n21081_o;
  wire n21083_o;
  wire n21085_o;
  wire n21087_o;
  wire n21089_o;
  wire n21091_o;
  wire n21093_o;
  wire n21095_o;
  wire n21097_o;
  wire n21099_o;
  wire n21101_o;
  wire n21103_o;
  wire n21105_o;
  wire n21107_o;
  wire n21109_o;
  wire n21111_o;
  wire n21113_o;
  wire n21115_o;
  wire [22:0] n21116_o;
  wire [22:0] n21129_o;
  wire [22:0] n21131_o;
  wire [22:0] n21133_o;
  wire [63:0] n21136_o;
  wire n21145_o;
  wire n21146_o;
  wire n21147_o;
  wire n21148_o;
  wire n21150_o;
  wire n21152_o;
  wire n21153_o;
  wire n21154_o;
  wire n21155_o;
  wire n21156_o;
  wire n21157_o;
  wire n21158_o;
  wire n21159_o;
  wire n21160_o;
  wire n21161_o;
  wire n21162_o;
  wire n21163_o;
  wire n21164_o;
  wire n21165_o;
  wire n21166_o;
  wire n21167_o;
  wire n21168_o;
  wire n21169_o;
  wire n21170_o;
  wire n21171_o;
  wire n21172_o;
  wire n21173_o;
  wire n21174_o;
  wire n21175_o;
  wire n21176_o;
  wire n21177_o;
  wire n21178_o;
  wire n21179_o;
  wire n21180_o;
  wire n21181_o;
  wire n21182_o;
  wire n21183_o;
  wire n21184_o;
  wire n21185_o;
  wire n21186_o;
  wire n21187_o;
  wire n21188_o;
  wire n21189_o;
  wire n21190_o;
  wire n21191_o;
  wire n21192_o;
  wire n21193_o;
  wire n21194_o;
  wire n21195_o;
  wire n21196_o;
  wire n21197_o;
  wire n21198_o;
  wire n21199_o;
  wire n21200_o;
  wire n21201_o;
  wire n21202_o;
  wire n21203_o;
  wire n21204_o;
  wire n21205_o;
  wire n21206_o;
  wire n21207_o;
  wire n21208_o;
  wire n21209_o;
  wire n21210_o;
  wire n21211_o;
  wire n21212_o;
  wire n21213_o;
  wire n21214_o;
  wire n21215_o;
  wire n21216_o;
  wire n21217_o;
  wire n21218_o;
  wire n21219_o;
  wire n21220_o;
  wire n21221_o;
  wire n21222_o;
  wire n21223_o;
  wire n21224_o;
  wire n21225_o;
  wire n21226_o;
  wire n21227_o;
  wire n21228_o;
  wire n21229_o;
  wire n21230_o;
  wire n21231_o;
  wire n21232_o;
  wire n21233_o;
  wire n21234_o;
  wire n21235_o;
  wire n21236_o;
  wire n21237_o;
  wire n21238_o;
  wire n21239_o;
  wire n21240_o;
  wire n21241_o;
  wire n21242_o;
  wire n21243_o;
  wire n21244_o;
  wire n21245_o;
  wire n21246_o;
  wire n21247_o;
  wire n21248_o;
  wire n21249_o;
  wire n21250_o;
  wire n21251_o;
  wire n21252_o;
  wire n21253_o;
  wire n21254_o;
  wire n21255_o;
  wire n21256_o;
  wire n21257_o;
  wire n21258_o;
  wire n21259_o;
  wire n21260_o;
  wire n21261_o;
  wire n21262_o;
  wire n21263_o;
  wire n21264_o;
  wire n21265_o;
  wire n21266_o;
  wire n21267_o;
  wire n21268_o;
  wire n21269_o;
  wire n21270_o;
  wire n21271_o;
  wire n21272_o;
  wire n21273_o;
  wire n21274_o;
  wire n21275_o;
  wire n21276_o;
  wire n21277_o;
  wire n21278_o;
  wire n21279_o;
  wire n21280_o;
  wire n21281_o;
  wire n21282_o;
  wire n21283_o;
  wire n21284_o;
  wire n21285_o;
  wire n21286_o;
  wire n21287_o;
  wire n21288_o;
  wire n21289_o;
  wire n21290_o;
  wire n21291_o;
  wire n21292_o;
  wire n21293_o;
  wire n21294_o;
  wire n21295_o;
  wire n21296_o;
  wire n21297_o;
  wire n21298_o;
  wire n21299_o;
  wire n21300_o;
  wire n21301_o;
  wire n21302_o;
  wire n21303_o;
  wire n21304_o;
  wire n21305_o;
  wire n21306_o;
  wire n21309_o;
  wire n21310_o;
  wire n21311_o;
  wire n21312_o;
  wire n21314_o;
  wire n21316_o;
  wire n21317_o;
  wire n21318_o;
  wire n21319_o;
  wire n21320_o;
  wire n21321_o;
  wire n21322_o;
  wire n21323_o;
  wire n21324_o;
  wire n21325_o;
  wire n21326_o;
  wire n21327_o;
  wire n21328_o;
  wire n21329_o;
  wire n21330_o;
  wire n21331_o;
  wire n21332_o;
  wire n21333_o;
  wire n21334_o;
  wire n21335_o;
  wire n21336_o;
  wire n21337_o;
  wire n21338_o;
  wire n21339_o;
  wire n21340_o;
  wire n21341_o;
  wire n21342_o;
  wire n21343_o;
  wire n21344_o;
  wire n21345_o;
  wire n21346_o;
  wire n21347_o;
  wire n21348_o;
  wire n21349_o;
  wire n21350_o;
  wire n21351_o;
  wire n21352_o;
  wire n21353_o;
  wire n21354_o;
  wire n21355_o;
  wire n21356_o;
  wire n21357_o;
  wire n21358_o;
  wire n21359_o;
  wire n21360_o;
  wire n21361_o;
  wire n21362_o;
  wire n21363_o;
  wire n21364_o;
  wire n21365_o;
  wire n21366_o;
  wire n21367_o;
  wire n21368_o;
  wire n21369_o;
  wire n21370_o;
  wire n21371_o;
  wire n21372_o;
  wire n21373_o;
  wire n21374_o;
  wire n21375_o;
  wire n21376_o;
  wire n21377_o;
  wire n21378_o;
  wire n21379_o;
  wire n21380_o;
  wire n21381_o;
  wire n21382_o;
  wire n21383_o;
  wire n21384_o;
  wire n21385_o;
  wire n21386_o;
  wire n21387_o;
  wire n21388_o;
  wire n21389_o;
  wire n21390_o;
  wire n21392_o;
  wire n21393_o;
  wire n21394_o;
  wire n21395_o;
  wire n21397_o;
  wire n21399_o;
  wire n21400_o;
  wire n21401_o;
  wire n21402_o;
  wire n21403_o;
  wire n21404_o;
  wire n21405_o;
  wire n21406_o;
  wire n21407_o;
  wire n21408_o;
  wire n21409_o;
  wire n21410_o;
  wire n21411_o;
  wire n21412_o;
  wire n21413_o;
  wire n21414_o;
  wire n21415_o;
  wire n21416_o;
  wire n21417_o;
  wire n21418_o;
  wire n21419_o;
  wire n21420_o;
  wire n21421_o;
  wire n21422_o;
  wire n21423_o;
  wire n21424_o;
  wire n21425_o;
  wire n21426_o;
  wire n21427_o;
  wire n21428_o;
  wire n21429_o;
  wire n21430_o;
  wire n21431_o;
  wire n21432_o;
  wire n21433_o;
  wire n21435_o;
  wire n21436_o;
  wire n21437_o;
  wire n21438_o;
  wire n21440_o;
  wire n21442_o;
  wire n21443_o;
  wire n21444_o;
  wire n21445_o;
  wire n21446_o;
  wire n21447_o;
  wire n21448_o;
  wire n21449_o;
  wire n21450_o;
  wire n21451_o;
  wire n21452_o;
  wire n21453_o;
  wire n21454_o;
  wire n21455_o;
  wire n21456_o;
  wire n21458_o;
  wire n21459_o;
  wire n21460_o;
  wire n21461_o;
  wire n21463_o;
  wire n21465_o;
  wire n21466_o;
  wire n21467_o;
  wire n21468_o;
  wire n21469_o;
  wire n21471_o;
  wire n21472_o;
  wire n21473_o;
  wire n21474_o;
  wire n21476_o;
  wire [5:0] n21478_o;
  wire [63:0] n21481_o;
  wire n21490_o;
  wire n21491_o;
  wire n21493_o;
  wire n21495_o;
  wire n21496_o;
  wire n21497_o;
  wire n21498_o;
  wire n21499_o;
  wire n21500_o;
  wire n21501_o;
  wire n21502_o;
  wire n21503_o;
  wire n21504_o;
  wire n21505_o;
  wire n21506_o;
  wire n21507_o;
  wire n21508_o;
  wire n21509_o;
  wire n21510_o;
  wire n21511_o;
  wire n21512_o;
  wire n21513_o;
  wire n21514_o;
  wire n21515_o;
  wire n21516_o;
  wire n21517_o;
  wire n21518_o;
  wire n21519_o;
  wire n21520_o;
  wire n21521_o;
  wire n21522_o;
  wire n21523_o;
  wire n21524_o;
  wire n21525_o;
  wire n21526_o;
  wire n21527_o;
  wire n21528_o;
  wire n21529_o;
  wire n21530_o;
  wire n21531_o;
  wire n21532_o;
  wire n21533_o;
  wire n21534_o;
  wire n21535_o;
  wire n21536_o;
  wire n21537_o;
  wire n21538_o;
  wire n21539_o;
  wire n21540_o;
  wire n21541_o;
  wire n21542_o;
  wire n21543_o;
  wire n21544_o;
  wire n21545_o;
  wire n21546_o;
  wire n21547_o;
  wire n21548_o;
  wire n21549_o;
  wire n21550_o;
  wire n21551_o;
  wire n21552_o;
  wire n21553_o;
  wire n21554_o;
  wire n21555_o;
  wire n21556_o;
  wire n21557_o;
  wire n21558_o;
  wire n21559_o;
  wire n21560_o;
  wire n21561_o;
  wire n21562_o;
  wire n21563_o;
  wire n21564_o;
  wire n21565_o;
  wire n21566_o;
  wire n21567_o;
  wire n21568_o;
  wire n21569_o;
  wire n21570_o;
  wire n21571_o;
  wire n21572_o;
  wire n21573_o;
  wire n21574_o;
  wire n21575_o;
  wire n21576_o;
  wire n21577_o;
  wire n21578_o;
  wire n21579_o;
  wire n21580_o;
  wire n21581_o;
  wire n21582_o;
  wire n21583_o;
  wire n21584_o;
  wire n21585_o;
  wire n21586_o;
  wire n21587_o;
  wire [1:0] n21590_o;
  wire n21591_o;
  wire n21593_o;
  wire [1:0] n21595_o;
  wire n21596_o;
  wire n21597_o;
  wire [1:0] n21598_o;
  wire n21599_o;
  wire n21600_o;
  wire [1:0] n21601_o;
  wire n21602_o;
  wire n21603_o;
  wire [1:0] n21604_o;
  wire n21605_o;
  wire n21606_o;
  wire [1:0] n21607_o;
  wire n21608_o;
  wire n21609_o;
  wire [1:0] n21610_o;
  wire n21611_o;
  wire n21612_o;
  wire [1:0] n21613_o;
  wire n21614_o;
  wire n21615_o;
  wire [1:0] n21616_o;
  wire n21617_o;
  wire n21618_o;
  wire [1:0] n21619_o;
  wire n21620_o;
  wire n21621_o;
  wire [1:0] n21622_o;
  wire n21623_o;
  wire n21624_o;
  wire [1:0] n21625_o;
  wire n21626_o;
  wire n21627_o;
  wire [1:0] n21628_o;
  wire n21629_o;
  wire n21630_o;
  wire [1:0] n21631_o;
  wire n21632_o;
  wire n21633_o;
  wire [1:0] n21634_o;
  wire n21635_o;
  wire n21636_o;
  wire [1:0] n21637_o;
  wire n21638_o;
  wire n21639_o;
  wire [3:0] n21641_o;
  wire n21642_o;
  wire n21644_o;
  wire [3:0] n21646_o;
  wire n21647_o;
  wire n21648_o;
  wire [3:0] n21649_o;
  wire n21650_o;
  wire n21651_o;
  wire [3:0] n21652_o;
  wire n21653_o;
  wire n21654_o;
  wire [3:0] n21655_o;
  wire n21656_o;
  wire n21657_o;
  wire [3:0] n21658_o;
  wire n21659_o;
  wire n21660_o;
  wire [3:0] n21661_o;
  wire n21662_o;
  wire n21663_o;
  wire [3:0] n21664_o;
  wire n21665_o;
  wire n21666_o;
  wire [7:0] n21668_o;
  wire n21669_o;
  wire n21671_o;
  wire [7:0] n21673_o;
  wire n21674_o;
  wire n21675_o;
  wire [7:0] n21676_o;
  wire n21677_o;
  wire n21678_o;
  wire [7:0] n21679_o;
  wire n21680_o;
  wire n21681_o;
  wire [15:0] n21683_o;
  wire n21684_o;
  wire n21686_o;
  wire [15:0] n21688_o;
  wire n21689_o;
  wire n21690_o;
  wire [31:0] n21692_o;
  wire n21693_o;
  wire n21695_o;
  wire [5:0] n21697_o;
  wire [3:0] n21699_o;
  wire [1:0] n21700_o;
  wire [5:0] n21701_o;
  wire n21704_o;
  wire [272:0] n21705_o;
  wire n21706_o;
  wire n21707_o;
  wire [63:0] n21708_o;
  wire [63:0] n21709_o;
  wire [63:0] n21710_o;
  wire [95:0] n21711_o;
  wire [272:0] n21712_o;
  wire n21713_o;
  wire [272:0] n21714_o;
  wire n21715_o;
  wire n21716_o;
  wire n21717_o;
  wire n21718_o;
  wire n21719_o;
  wire n21720_o;
  wire n21721_o;
  wire n21722_o;
  wire [31:0] n21723_o;
  wire [63:0] n21725_o;
  wire [63:0] n21726_o;
  wire [63:0] n21727_o;
  wire [63:0] n21728_o;
  wire [63:0] n21729_o;
  wire n21732_o;
  wire [63:0] n21734_o;
  wire [272:0] n21735_o;
  wire n21736_o;
  wire n21739_o;
  wire [272:0] n21740_o;
  wire n21741_o;
  wire n21743_o;
  wire [272:0] n21744_o;
  wire n21745_o;
  wire n21748_o;
  wire n21750_o;
  wire n21753_o;
  wire n21756_o;
  wire [63:0] n21759_o;
  wire [1:0] n21761_o;
  wire n21762_o;
  wire [272:0] n21763_o;
  wire n21764_o;
  wire n21765_o;
  wire [272:0] n21766_o;
  wire n21767_o;
  wire n21768_o;
  wire [272:0] n21769_o;
  wire n21770_o;
  wire [272:0] n21771_o;
  wire n21772_o;
  wire n21773_o;
  wire n21774_o;
  wire [272:0] n21775_o;
  wire n21776_o;
  wire n21778_o;
  wire [272:0] n21781_o;
  wire n21782_o;
  wire [272:0] n21783_o;
  wire n21784_o;
  wire n21785_o;
  wire [1:0] n21786_o;
  wire [1:0] n21787_o;
  wire n21788_o;
  wire n21789_o;
  wire n21791_o;
  wire n21792_o;
  wire n21793_o;
  wire n21794_o;
  wire n21797_o;
  wire n21799_o;
  wire n21800_o;
  wire n21801_o;
  wire n21802_o;
  wire n21804_o;
  wire n21805_o;
  wire n21806_o;
  wire [272:0] n21807_o;
  wire n21808_o;
  wire n21809_o;
  wire n21810_o;
  wire [1:0] n21813_o;
  wire n21814_o;
  wire n21815_o;
  wire n21818_o;
  wire n21820_o;
  wire n21822_o;
  wire n21824_o;
  wire [1:0] n21825_o;
  wire n21826_o;
  wire n21827_o;
  wire n21829_o;
  wire n21830_o;
  wire n21832_o;
  wire n21834_o;
  wire [272:0] n21835_o;
  wire n21836_o;
  wire [272:0] n21837_o;
  wire n21838_o;
  wire [272:0] n21839_o;
  wire n21840_o;
  wire n21841_o;
  wire [272:0] n21842_o;
  wire n21843_o;
  wire [272:0] n21844_o;
  wire n21845_o;
  wire [1:0] n21849_o;
  wire n21850_o;
  wire n21851_o;
  wire [272:0] n21852_o;
  wire n21853_o;
  wire n21854_o;
  wire n21855_o;
  wire [31:0] n21856_o;
  wire [272:0] n21857_o;
  wire [63:0] n21858_o;
  wire [63:0] n21859_o;
  wire [63:0] n21860_o;
  wire [31:0] n21861_o;
  wire [31:0] n21862_o;
  wire [95:0] n21863_o;
  wire [95:0] n21864_o;
  wire [1:0] n21865_o;
  wire [95:0] n21866_o;
  wire n21868_o;
  wire n21869_o;
  wire n21871_o;
  wire n21872_o;
  wire [95:0] n21873_o;
  wire n21875_o;
  wire n21876_o;
  wire n21878_o;
  wire n21880_o;
  wire n21881_o;
  wire [272:0] n21882_o;
  wire n21883_o;
  wire n21884_o;
  wire [1:0] n21887_o;
  wire [1:0] n21888_o;
  wire n21889_o;
  wire n21890_o;
  wire n21893_o;
  wire n21895_o;
  wire n21897_o;
  wire n21899_o;
  wire n21900_o;
  wire n21901_o;
  wire n21902_o;
  wire [272:0] n21903_o;
  wire n21904_o;
  wire [272:0] n21905_o;
  wire n21906_o;
  wire n21907_o;
  wire n21908_o;
  wire n21909_o;
  wire n21911_o;
  wire [1:0] n21912_o;
  wire [1:0] n21914_o;
  wire n21916_o;
  wire n21918_o;
  wire n21920_o;
  wire n21922_o;
  wire n21924_o;
  wire n21926_o;
  wire [3:0] n21927_o;
  wire [1:0] n21928_o;
  reg [1:0] n21930_o;
  reg n21932_o;
  reg [95:0] n21934_o;
  wire n21935_o;
  reg n21937_o;
  wire n21938_o;
  reg n21940_o;
  wire [81:0] n21941_o;
  reg n21946_o;
  reg n21950_o;
  reg n21954_o;
  reg n21958_o;
  reg n21960_o;
  reg n21963_o;
  reg n21966_o;
  reg [1:0] n21969_o;
  reg n21972_o;
  reg n21975_o;
  reg n21978_o;
  reg n21981_o;
  localparam [31:0] n21982_o = 32'b00000000000000000000000000000000;
  wire [17:0] n21984_o;
  wire [4:0] n21986_o;
  wire n21988_o;
  wire n21990_o;
  wire n21991_o;
  wire n21992_o;
  wire [1:0] n21995_o;
  wire n21996_o;
  wire [272:0] n21997_o;
  wire n21998_o;
  wire n21999_o;
  wire [272:0] n22001_o;
  wire n22002_o;
  wire [272:0] n22003_o;
  wire n22004_o;
  wire n22005_o;
  wire n22006_o;
  wire [75:0] n22007_o;
  wire [272:0] n22008_o;
  wire [63:0] n22009_o;
  wire [272:0] n22010_o;
  wire n22011_o;
  wire [272:0] n22013_o;
  wire [63:0] n22014_o;
  wire [272:0] n22015_o;
  wire n22016_o;
  wire n22017_o;
  wire [272:0] n22018_o;
  wire [63:0] n22019_o;
  wire n22020_o;
  wire n22021_o;
  wire [31:0] n22023_o;
  wire [31:0] n22025_o;
  wire [31:0] n22026_o;
  wire [11:0] n22027_o;
  wire n22028_o;
  wire n22029_o;
  wire n22030_o;
  wire n22031_o;
  wire n22032_o;
  wire n22033_o;
  wire [1:0] n22036_o;
  wire [11:0] n22037_o;
  wire [1:0] n22038_o;
  wire [1:0] n22039_o;
  wire n22040_o;
  wire n22041_o;
  wire n22042_o;
  wire n22043_o;
  wire [95:0] n22044_o;
  wire [95:0] n22045_o;
  wire [11:0] n22046_o;
  wire [1:0] n22047_o;
  wire [1:0] n22048_o;
  wire n22049_o;
  wire n22050_o;
  wire n22051_o;
  wire n22052_o;
  wire [63:0] n22053_o;
  wire [63:0] n22054_o;
  wire [31:0] n22055_o;
  wire [31:0] n22056_o;
  wire [31:0] n22057_o;
  wire [11:0] n22058_o;
  wire [1:0] n22059_o;
  wire [1:0] n22060_o;
  wire n22061_o;
  wire n22062_o;
  wire n22063_o;
  wire n22064_o;
  wire [95:0] n22065_o;
  wire [75:0] n22066_o;
  wire [95:0] n22067_o;
  wire [75:0] n22068_o;
  wire [1:0] n22069_o;
  wire [1:0] n22070_o;
  wire n22071_o;
  wire n22072_o;
  wire n22073_o;
  wire n22074_o;
  wire [1:0] n22076_o;
  wire [7:0] n22078_o;
  wire n22079_o;
  wire n22080_o;
  wire [1:0] n22081_o;
  wire n22083_o;
  wire [63:0] n22084_o;
  wire n22086_o;
  wire n22088_o;
  wire [63:0] n22089_o;
  wire [2:0] n22090_o;
  reg [63:0] n22091_o;
  wire n22092_o;
  wire n22093_o;
  wire n22094_o;
  wire n22095_o;
  wire n22096_o;
  wire n22097_o;
  wire [63:0] n22098_o;
  wire [7:0] n22099_o;
  wire n22100_o;
  wire n22101_o;
  wire [272:0] n22102_o;
  wire n22103_o;
  wire [272:0] n22104_o;
  wire n22105_o;
  wire [272:0] n22106_o;
  wire n22107_o;
  wire [272:0] n22108_o;
  wire n22109_o;
  wire [272:0] n22110_o;
  wire n22111_o;
  wire [272:0] n22112_o;
  wire n22113_o;
  wire [272:0] n22114_o;
  wire [63:0] n22115_o;
  wire [272:0] n22116_o;
  wire [7:0] n22117_o;
  wire [272:0] n22118_o;
  wire n22119_o;
  wire [272:0] n22120_o;
  wire n22121_o;
  wire [71:0] n22122_o;
  wire [71:0] n22123_o;
  wire n22124_o;
  wire [71:0] n22125_o;
  wire [7:0] n22126_o;
  wire [272:0] n22127_o;
  wire [63:0] n22128_o;
  wire [63:0] n22129_o;
  wire [272:0] n22130_o;
  wire n22131_o;
  wire [272:0] n22132_o;
  wire n22133_o;
  wire n22134_o;
  wire n22135_o;
  wire n22136_o;
  wire [272:0] n22137_o;
  wire n22138_o;
  wire [272:0] n22139_o;
  wire n22140_o;
  wire [272:0] n22141_o;
  wire n22142_o;
  wire [272:0] n22143_o;
  wire n22144_o;
  wire [272:0] n22145_o;
  wire [9:0] n22146_o;
  wire [272:0] n22147_o;
  wire [63:0] n22148_o;
  wire [272:0] n22149_o;
  wire n22150_o;
  wire [272:0] n22151_o;
  wire [63:0] n22152_o;
  wire [272:0] n22153_o;
  wire [2:0] n22154_o;
  wire n22155_o;
  wire [272:0] n22156_o;
  wire [6:0] n22157_o;
  wire [272:0] n22158_o;
  wire [4:0] n22159_o;
  wire [272:0] n22160_o;
  wire n22161_o;
  wire n22162_o;
  wire n22163_o;
  wire n22164_o;
  wire [11:0] n22165_o;
  wire [63:0] n22166_o;
  wire [15:0] n22167_o;
  wire n22168_o;
  wire [2:0] n22169_o;
  wire [272:0] n22170_o;
  wire n22171_o;
  wire n22172_o;
  wire n22173_o;
  wire n22174_o;
  wire n22175_o;
  wire [380:0] n22176_o;
  reg [337:0] n22184_q;
  reg [373:0] n22185_q;
  reg [380:0] n22186_q;
  reg n22187_q;
  wire [31:0] n22188_o;
  wire [63:0] n22189_o;
  wire [63:0] n22190_o;
  reg n22191_q;
  wire [2:0] n22192_o;
  wire [175:0] n22193_o;
  wire [145:0] n22194_o;
  wire [144:0] n22195_o;
  localparam [9:0] n22196_o = 10'bZ;
  wire [7:0] n22197_o;
  wire [7:0] n22198_o;
  wire [7:0] n22199_o;
  wire [7:0] n22200_o;
  wire [7:0] n22201_o;
  wire [7:0] n22202_o;
  wire [7:0] n22203_o;
  wire [7:0] n22204_o;
  wire [1:0] n22205_o;
  reg [7:0] n22206_o;
  wire [1:0] n22207_o;
  reg [7:0] n22208_o;
  wire n22209_o;
  wire [7:0] n22210_o;
  wire [7:0] n22211_o;
  wire [7:0] n22212_o;
  wire [7:0] n22213_o;
  wire [7:0] n22214_o;
  wire [7:0] n22215_o;
  wire [7:0] n22216_o;
  wire [7:0] n22217_o;
  wire [7:0] n22218_o;
  wire [1:0] n22219_o;
  reg [7:0] n22220_o;
  wire [1:0] n22221_o;
  reg [7:0] n22222_o;
  wire n22223_o;
  wire [7:0] n22224_o;
  wire [7:0] n22225_o;
  wire [7:0] n22226_o;
  wire [7:0] n22227_o;
  wire [7:0] n22228_o;
  wire [7:0] n22229_o;
  wire [7:0] n22230_o;
  wire [7:0] n22231_o;
  wire [7:0] n22232_o;
  wire [1:0] n22233_o;
  reg [7:0] n22234_o;
  wire [1:0] n22235_o;
  reg [7:0] n22236_o;
  wire n22237_o;
  wire [7:0] n22238_o;
  wire [7:0] n22239_o;
  wire [7:0] n22240_o;
  wire [7:0] n22241_o;
  wire [7:0] n22242_o;
  wire [7:0] n22243_o;
  wire [7:0] n22244_o;
  wire [7:0] n22245_o;
  wire [7:0] n22246_o;
  wire [1:0] n22247_o;
  reg [7:0] n22248_o;
  wire [1:0] n22249_o;
  reg [7:0] n22250_o;
  wire n22251_o;
  wire [7:0] n22252_o;
  wire [7:0] n22253_o;
  wire [7:0] n22254_o;
  wire [7:0] n22255_o;
  wire [7:0] n22256_o;
  wire [7:0] n22257_o;
  wire [7:0] n22258_o;
  wire [7:0] n22259_o;
  wire [7:0] n22260_o;
  wire [1:0] n22261_o;
  reg [7:0] n22262_o;
  wire [1:0] n22263_o;
  reg [7:0] n22264_o;
  wire n22265_o;
  wire [7:0] n22266_o;
  wire [7:0] n22267_o;
  wire [7:0] n22268_o;
  wire [7:0] n22269_o;
  wire [7:0] n22270_o;
  wire [7:0] n22271_o;
  wire [7:0] n22272_o;
  wire [7:0] n22273_o;
  wire [7:0] n22274_o;
  wire [1:0] n22275_o;
  reg [7:0] n22276_o;
  wire [1:0] n22277_o;
  reg [7:0] n22278_o;
  wire n22279_o;
  wire [7:0] n22280_o;
  wire [7:0] n22281_o;
  wire [7:0] n22282_o;
  wire [7:0] n22283_o;
  wire [7:0] n22284_o;
  wire [7:0] n22285_o;
  wire [7:0] n22286_o;
  wire [7:0] n22287_o;
  wire [7:0] n22288_o;
  wire [1:0] n22289_o;
  reg [7:0] n22290_o;
  wire [1:0] n22291_o;
  reg [7:0] n22292_o;
  wire n22293_o;
  wire [7:0] n22294_o;
  wire [7:0] n22295_o;
  wire [7:0] n22296_o;
  wire [7:0] n22297_o;
  wire [7:0] n22298_o;
  wire [7:0] n22299_o;
  wire [7:0] n22300_o;
  wire [7:0] n22301_o;
  wire [7:0] n22302_o;
  wire [1:0] n22303_o;
  reg [7:0] n22304_o;
  wire [1:0] n22305_o;
  reg [7:0] n22306_o;
  wire n22307_o;
  wire [7:0] n22308_o;
  wire [7:0] n22309_o;
  wire [7:0] n22310_o;
  wire [7:0] n22311_o;
  wire [7:0] n22312_o;
  wire [7:0] n22313_o;
  wire [7:0] n22314_o;
  wire [7:0] n22315_o;
  wire [7:0] n22316_o;
  wire [1:0] n22317_o;
  reg [7:0] n22318_o;
  wire [1:0] n22319_o;
  reg [7:0] n22320_o;
  wire n22321_o;
  wire [7:0] n22322_o;
  wire [7:0] n22323_o;
  wire [7:0] n22324_o;
  wire [7:0] n22325_o;
  wire [7:0] n22326_o;
  wire [7:0] n22327_o;
  wire [7:0] n22328_o;
  wire [7:0] n22329_o;
  wire [7:0] n22330_o;
  wire [1:0] n22331_o;
  reg [7:0] n22332_o;
  wire [1:0] n22333_o;
  reg [7:0] n22334_o;
  wire n22335_o;
  wire [7:0] n22336_o;
  wire [7:0] n22337_o;
  wire [7:0] n22338_o;
  wire [7:0] n22339_o;
  wire [7:0] n22340_o;
  wire [7:0] n22341_o;
  wire [7:0] n22342_o;
  wire [7:0] n22343_o;
  wire [7:0] n22344_o;
  wire [1:0] n22345_o;
  reg [7:0] n22346_o;
  wire [1:0] n22347_o;
  reg [7:0] n22348_o;
  wire n22349_o;
  wire [7:0] n22350_o;
  wire [7:0] n22351_o;
  wire [7:0] n22352_o;
  wire [7:0] n22353_o;
  wire [7:0] n22354_o;
  wire [7:0] n22355_o;
  wire [7:0] n22356_o;
  wire [7:0] n22357_o;
  wire [7:0] n22358_o;
  wire [1:0] n22359_o;
  reg [7:0] n22360_o;
  wire [1:0] n22361_o;
  reg [7:0] n22362_o;
  wire n22363_o;
  wire [7:0] n22364_o;
  wire [7:0] n22365_o;
  wire [7:0] n22366_o;
  wire [7:0] n22367_o;
  wire [7:0] n22368_o;
  wire [7:0] n22369_o;
  wire [7:0] n22370_o;
  wire [7:0] n22371_o;
  wire [7:0] n22372_o;
  wire [1:0] n22373_o;
  reg [7:0] n22374_o;
  wire [1:0] n22375_o;
  reg [7:0] n22376_o;
  wire n22377_o;
  wire [7:0] n22378_o;
  wire [7:0] n22379_o;
  wire [7:0] n22380_o;
  wire [7:0] n22381_o;
  wire [7:0] n22382_o;
  wire [7:0] n22383_o;
  wire [7:0] n22384_o;
  wire [7:0] n22385_o;
  wire [7:0] n22386_o;
  wire [1:0] n22387_o;
  reg [7:0] n22388_o;
  wire [1:0] n22389_o;
  reg [7:0] n22390_o;
  wire n22391_o;
  wire [7:0] n22392_o;
  wire [7:0] n22393_o;
  wire [7:0] n22394_o;
  wire [7:0] n22395_o;
  wire [7:0] n22396_o;
  wire [7:0] n22397_o;
  wire [7:0] n22398_o;
  wire [7:0] n22399_o;
  wire [7:0] n22400_o;
  wire [1:0] n22401_o;
  reg [7:0] n22402_o;
  wire [1:0] n22403_o;
  reg [7:0] n22404_o;
  wire n22405_o;
  wire [7:0] n22406_o;
  wire [7:0] n22407_o;
  wire [7:0] n22408_o;
  wire [7:0] n22409_o;
  wire [7:0] n22410_o;
  wire [7:0] n22411_o;
  wire [7:0] n22412_o;
  wire [7:0] n22413_o;
  wire [7:0] n22414_o;
  wire [1:0] n22415_o;
  reg [7:0] n22416_o;
  wire [1:0] n22417_o;
  reg [7:0] n22418_o;
  wire n22419_o;
  wire [7:0] n22420_o;
  assign e_out_busy = n19328_o;
  assign e_out_in_progress = n19329_o;
  assign e_out_interrupt = n19330_o;
  assign l_out_valid = n19332_o;
  assign l_out_instr_tag = n19333_o;
  assign l_out_write_enable = n19334_o;
  assign l_out_write_reg = n19335_o;
  assign l_out_write_data = n19336_o;
  assign l_out_xerc = n19337_o;
  assign l_out_rc = n19338_o;
  assign l_out_store_done = n19339_o;
  assign l_out_interrupt = n19340_o;
  assign l_out_intr_vec = n19341_o;
  assign l_out_srr0 = n19342_o;
  assign l_out_srr1 = n19343_o;
  assign d_out_valid = n19345_o;
  assign d_out_hold = n19346_o;
  assign d_out_load = n19347_o;
  assign d_out_dcbz = n19348_o;
  assign d_out_nc = n19349_o;
  assign d_out_reserve = n19350_o;
  assign d_out_atomic = n19351_o;
  assign d_out_atomic_last = n19352_o;
  assign d_out_virt_mode = n19353_o;
  assign d_out_priv_mode = n19354_o;
  assign d_out_addr = n19355_o;
  assign d_out_data = n19356_o;
  assign d_out_byte_sel = n19357_o;
  assign m_out_valid = n19360_o;
  assign m_out_tlbie = n19361_o;
  assign m_out_slbia = n19362_o;
  assign m_out_mtspr = n19363_o;
  assign m_out_iside = n19364_o;
  assign m_out_load = n19365_o;
  assign m_out_priv = n19366_o;
  assign m_out_sprn = n19367_o;
  assign m_out_addr = n19368_o;
  assign m_out_rs = n19369_o;
  assign events_load_complete = n19372_o;
  assign events_store_complete = n19373_o;
  assign events_itlb_miss = n19374_o;
  assign log_out = n22196_o;
  assign n19326_o = {l_in_msr, l_in_second, l_in_repeat, l_in_is_32bit, l_in_mode_32bit, l_in_priv_mode, l_in_virt_mode, l_in_rc, l_in_reserve, l_in_xerc, l_in_update, l_in_sign_extend, l_in_byte_reverse, l_in_ci, l_in_length, l_in_write_reg, l_in_data, l_in_addr2, l_in_addr1, l_in_instr_tag, l_in_insn, l_in_nia, l_in_op, l_in_valid};
  /* fpu.vhdl:22:9  */
  assign n19328_o = n22192_o[0];
  /* fpu.vhdl:20:9  */
  assign n19329_o = n22192_o[1];
  /* fpu.vhdl:544:9  */
  assign n19330_o = n22192_o[2];
  assign n19332_o = n22193_o[0];
  assign n19333_o = n22193_o[3:1];
  assign n19334_o = n22193_o[4];
  assign n19335_o = n22193_o[11:5];
  /* fpu.vhdl:519:14  */
  assign n19336_o = n22193_o[75:12];
  /* fpu.vhdl:519:14  */
  assign n19337_o = n22193_o[80:76];
  assign n19338_o = n22193_o[81];
  /* fpu.vhdl:519:14  */
  assign n19339_o = n22193_o[82];
  assign n19340_o = n22193_o[83];
  assign n19341_o = n22193_o[95:84];
  assign n19342_o = n22193_o[159:96];
  assign n19343_o = n22193_o[175:160];
  assign n19345_o = n22194_o[0];
  /* fpu.vhdl:449:14  */
  assign n19346_o = n22194_o[1];
  /* fpu.vhdl:449:14  */
  assign n19347_o = n22194_o[2];
  assign n19348_o = n22194_o[3];
  /* fpu.vhdl:449:14  */
  assign n19349_o = n22194_o[4];
  /* fpu.vhdl:2520:9  */
  assign n19350_o = n22194_o[5];
  assign n19351_o = n22194_o[6];
  assign n19352_o = n22194_o[7];
  assign n19353_o = n22194_o[8];
  assign n19354_o = n22194_o[9];
  assign n19355_o = n22194_o[73:10];
  assign n19356_o = n22194_o[137:74];
  assign n19357_o = n22194_o[145:138];
  /* loadstore1.vhdl:685:63  */
  assign n19358_o = {d_in_cache_paradox, d_in_error, d_in_store_done, d_in_data, d_in_valid};
  assign n19360_o = n22195_o[0];
  assign n19361_o = n22195_o[1];
  assign n19362_o = n22195_o[2];
  assign n19363_o = n22195_o[3];
  assign n19364_o = n22195_o[4];
  assign n19365_o = n22195_o[5];
  /* helpers.vhdl:237:18  */
  assign n19366_o = n22195_o[6];
  assign n19367_o = n22195_o[16:7];
  /* helpers.vhdl:236:18  */
  assign n19368_o = n22195_o[80:17];
  assign n19369_o = n22195_o[144:81];
  /* helpers.vhdl:235:18  */
  assign n19370_o = {m_in_sprval, m_in_rc_error, m_in_perm_error, m_in_segerr, m_in_badtree, m_in_invalid, m_in_err, m_in_done};
  /* helpers.vhdl:234:18  */
  assign n19372_o = n22169_o[0];
  assign n19373_o = n22169_o[1];
  /* helpers.vhdl:30:14  */
  assign n19374_o = n22169_o[2];
  /* loadstore1.vhdl:155:12  */
  assign req_in = n19943_o; // (signal)
  /* loadstore1.vhdl:156:12  */
  assign r1 = n22184_q; // (signal)
  /* loadstore1.vhdl:156:16  */
  assign r1in = n20166_o; // (signal)
  /* loadstore1.vhdl:157:12  */
  assign r2 = n22185_q; // (signal)
  /* loadstore1.vhdl:157:16  */
  assign r2in = n20475_o; // (signal)
  /* loadstore1.vhdl:158:12  */
  assign r3 = n22186_q; // (signal)
  /* loadstore1.vhdl:158:16  */
  assign r3in = n22176_o; // (signal)
  /* loadstore1.vhdl:160:12  */
  assign busy = n19970_o; // (signal)
  /* loadstore1.vhdl:161:12  */
  assign complete = n19981_o; // (signal)
  /* loadstore1.vhdl:162:12  */
  assign in_progress = n19988_o; // (signal)
  /* loadstore1.vhdl:163:12  */
  assign flushing = n22187_q; // (signal)
  /* loadstore1.vhdl:165:12  */
  assign store_sp_data = n22188_o; // (signal)
  /* loadstore1.vhdl:166:12  */
  assign load_dp_data = n22189_o; // (signal)
  /* loadstore1.vhdl:167:12  */
  assign store_data = n22190_o; // (signal)
  /* loadstore1.vhdl:169:12  */
  assign stage1_issue_enable = n20003_o; // (signal)
  /* loadstore1.vhdl:170:12  */
  assign stage1_req = n20165_o; // (signal)
  /* loadstore1.vhdl:171:12  */
  assign stage1_dcreq = n20163_o; // (signal)
  /* loadstore1.vhdl:172:12  */
  assign stage1_dreq = n22191_q; // (signal)
  /* loadstore1.vhdl:173:12  */
  assign stage2_busy_next = n20471_o; // (signal)
  /* loadstore1.vhdl:174:12  */
  assign stage3_busy_next = n22175_o; // (signal)
  /* loadstore1.vhdl:294:48  */
  assign n19390_o = r1in[272:0];
  /* loadstore1.vhdl:294:52  */
  assign n19391_o = n19390_o[0];
  /* loadstore1.vhdl:294:67  */
  assign n19392_o = r1in[272:0];
  /* loadstore1.vhdl:294:71  */
  assign n19393_o = n19392_o[206];
  /* loadstore1.vhdl:294:58  */
  assign n19394_o = n19391_o & n19393_o;
  /* loadstore1.vhdl:294:39  */
  assign n19395_o = flushing | n19394_o;
  /* loadstore1.vhdl:295:38  */
  assign n19396_o = r3in[285];
  /* loadstore1.vhdl:295:29  */
  assign n19397_o = ~n19396_o;
  /* loadstore1.vhdl:294:84  */
  assign n19398_o = n19395_o & n19397_o;
  /* helpers.vhdl:33:14  */
  assign n19399_o = r1in[0];
  /* loadstore1.vhdl:276:13  */
  assign n19400_o = rst ? 1'b0 : n19399_o;
  /* helpers.vhdl:33:14  */
  assign n19401_o = r1in[337:1];
  assign n19402_o = r1[337:1];
  /* loadstore1.vhdl:276:13  */
  assign n19403_o = rst ? n19402_o : n19401_o;
  assign n19404_o = {1'b0, 1'b0, 1'b0};
  assign n19405_o = r2in[0];
  /* loadstore1.vhdl:276:13  */
  assign n19406_o = rst ? 1'b0 : n19405_o;
  assign n19407_o = r2in[304:1];
  assign n19408_o = r2[304:1];
  /* loadstore1.vhdl:276:13  */
  assign n19409_o = rst ? n19408_o : n19407_o;
  assign n19410_o = r2in[307:305];
  /* loadstore1.vhdl:276:13  */
  assign n19411_o = rst ? n19404_o : n19410_o;
  assign n19412_o = r2in[373:308];
  assign n19413_o = r2[373:308];
  /* loadstore1.vhdl:276:13  */
  assign n19414_o = rst ? n19413_o : n19412_o;
  assign n19415_o = {32'b00000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000};
  assign n19416_o = {1'b0, 1'b1};
  assign n19417_o = r3in[1:0];
  /* loadstore1.vhdl:276:13  */
  assign n19418_o = rst ? 2'b00 : n19417_o;
  assign n19419_o = r3in[4:2];
  assign n19420_o = r3[4:2];
  /* loadstore1.vhdl:276:13  */
  assign n19421_o = rst ? n19420_o : n19419_o;
  assign n19422_o = r3in[5];
  /* loadstore1.vhdl:276:13  */
  assign n19423_o = rst ? 1'b0 : n19422_o;
  assign n19424_o = r3in[83:6];
  assign n19425_o = r3[83:6];
  /* loadstore1.vhdl:276:13  */
  assign n19426_o = rst ? n19425_o : n19424_o;
  assign n19427_o = r3in[84];
  /* loadstore1.vhdl:276:13  */
  assign n19428_o = rst ? 1'b0 : n19427_o;
  assign n19429_o = r3in[148:85];
  assign n19430_o = r3[148:85];
  /* loadstore1.vhdl:276:13  */
  assign n19431_o = rst ? n19430_o : n19429_o;
  assign n19432_o = r3in[244:149];
  /* loadstore1.vhdl:276:13  */
  assign n19433_o = rst ? n19415_o : n19432_o;
  assign n19434_o = r3in[283:245];
  assign n19435_o = r3[283:245];
  /* loadstore1.vhdl:276:13  */
  assign n19436_o = rst ? n19435_o : n19434_o;
  assign n19437_o = r3in[285:284];
  /* loadstore1.vhdl:276:13  */
  assign n19438_o = rst ? n19416_o : n19437_o;
  assign n19439_o = r3in[380:286];
  assign n19440_o = r3[380:286];
  /* loadstore1.vhdl:276:13  */
  assign n19441_o = rst ? n19440_o : n19439_o;
  /* loadstore1.vhdl:276:13  */
  assign n19443_o = rst ? 1'b0 : n19398_o;
  assign n19449_o = {n19403_o, n19400_o};
  assign n19451_o = {n19414_o, n19411_o, n19409_o, n19406_o};
  assign n19453_o = {n19441_o, n19438_o, n19436_o, n19433_o, n19431_o, n19428_o, n19426_o, n19423_o, n19421_o, n19418_o};
  /* loadstore1.vhdl:317:43  */
  assign n19462_o = n19326_o[297];
  /* loadstore1.vhdl:319:38  */
  assign n19464_o = n19326_o[296:286];
  /* loadstore1.vhdl:320:20  */
  assign n19466_o = $unsigned(n19464_o) > $unsigned(11'b01110000000);
  /* loadstore1.vhdl:321:47  */
  assign n19467_o = n19326_o[296];
  /* loadstore1.vhdl:322:56  */
  assign n19468_o = n19326_o[292:263];
  /* loadstore1.vhdl:323:23  */
  assign n19470_o = $unsigned(n19464_o) >= $unsigned(11'b01101101010);
  /* loadstore1.vhdl:325:40  */
  assign n19471_o = n19326_o[285:264];
  /* loadstore1.vhdl:325:29  */
  assign n19473_o = {1'b1, n19471_o};
  /* loadstore1.vhdl:326:33  */
  assign n19474_o = n19464_o[4:0];
  /* loadstore1.vhdl:326:28  */
  assign n19476_o = 5'b00000 - n19474_o;
  /* loadstore1.vhdl:212:19  */
  assign n19484_o = n19476_o[1:0];
  /* loadstore1.vhdl:213:13  */
  assign n19486_o = n19484_o == 2'b00;
  /* loadstore1.vhdl:216:34  */
  assign n19487_o = n19473_o[22:1];
  /* loadstore1.vhdl:216:28  */
  assign n19489_o = {1'b0, n19487_o};
  /* loadstore1.vhdl:215:13  */
  assign n19491_o = n19484_o == 2'b01;
  /* loadstore1.vhdl:218:35  */
  assign n19492_o = n19473_o[22:2];
  /* loadstore1.vhdl:218:29  */
  assign n19494_o = {2'b00, n19492_o};
  /* loadstore1.vhdl:217:13  */
  assign n19496_o = n19484_o == 2'b10;
  /* loadstore1.vhdl:220:36  */
  assign n19497_o = n19473_o[22:3];
  /* loadstore1.vhdl:220:30  */
  assign n19499_o = {3'b000, n19497_o};
  assign n19500_o = {n19496_o, n19491_o, n19486_o};
  /* loadstore1.vhdl:212:9  */
  always @*
    case (n19500_o)
      3'b100: n19501_o = n19494_o;
      3'b010: n19501_o = n19489_o;
      3'b001: n19501_o = n19473_o;
      default: n19501_o = n19499_o;
    endcase
  /* loadstore1.vhdl:222:19  */
  assign n19503_o = n19476_o[4:2];
  /* loadstore1.vhdl:223:13  */
  assign n19505_o = n19503_o == 3'b000;
  /* loadstore1.vhdl:226:34  */
  assign n19506_o = n19501_o[22:4];
  /* loadstore1.vhdl:226:29  */
  assign n19508_o = {4'b0000, n19506_o};
  /* loadstore1.vhdl:225:13  */
  assign n19510_o = n19503_o == 3'b001;
  /* loadstore1.vhdl:228:35  */
  assign n19511_o = n19501_o[22:8];
  /* loadstore1.vhdl:228:30  */
  assign n19513_o = {8'b00000000, n19511_o};
  /* loadstore1.vhdl:227:13  */
  assign n19515_o = n19503_o == 3'b010;
  /* loadstore1.vhdl:230:36  */
  assign n19516_o = n19501_o[22:12];
  /* loadstore1.vhdl:230:31  */
  assign n19518_o = {12'b000000000000, n19516_o};
  /* loadstore1.vhdl:229:13  */
  assign n19520_o = n19503_o == 3'b011;
  /* loadstore1.vhdl:232:37  */
  assign n19521_o = n19501_o[22:16];
  /* loadstore1.vhdl:232:32  */
  assign n19523_o = {16'b0000000000000000, n19521_o};
  /* loadstore1.vhdl:231:13  */
  assign n19525_o = n19503_o == 3'b100;
  /* loadstore1.vhdl:234:38  */
  assign n19526_o = n19501_o[22:20];
  /* loadstore1.vhdl:234:33  */
  assign n19528_o = {20'b00000000000000000000, n19526_o};
  assign n19529_o = {n19525_o, n19520_o, n19515_o, n19510_o, n19505_o};
  /* loadstore1.vhdl:222:9  */
  always @*
    case (n19529_o)
      5'b10000: n19530_o = n19523_o;
      5'b01000: n19530_o = n19518_o;
      5'b00100: n19530_o = n19513_o;
      5'b00010: n19530_o = n19508_o;
      5'b00001: n19530_o = n19501_o;
      default: n19530_o = n19528_o;
    endcase
  assign n19532_o = n19463_o[22:0];
  /* loadstore1.vhdl:323:13  */
  assign n19533_o = n19470_o ? n19530_o : n19532_o;
  assign n19536_o = {n19467_o, n19468_o};
  assign n19537_o = n19536_o[22:0];
  /* loadstore1.vhdl:320:13  */
  assign n19538_o = n19466_o ? n19537_o : n19533_o;
  assign n19539_o = n19536_o[30:23];
  assign n19540_o = n19463_o[30:23];
  /* loadstore1.vhdl:320:13  */
  assign n19541_o = n19466_o ? n19539_o : n19540_o;
  /* loadstore1.vhdl:340:34  */
  assign n19555_o = r3[267:245];
  /* loadstore1.vhdl:341:42  */
  assign n19556_o = r3[275:268];
  /* loadstore1.vhdl:342:40  */
  assign n19557_o = r3[275:268];
  /* loadstore1.vhdl:342:23  */
  assign n19558_o = |(n19557_o);
  /* loadstore1.vhdl:343:41  */
  assign n19559_o = r3[275:268];
  /* loadstore1.vhdl:343:23  */
  assign n19560_o = &(n19559_o);
  /* loadstore1.vhdl:348:33  */
  assign n19561_o = {3'b0, n19556_o};  //  uext
  /* loadstore1.vhdl:348:31  */
  assign n19563_o = 11'b01110000000 + n19561_o;
  /* loadstore1.vhdl:349:22  */
  assign n19564_o = r3[277];
  /* loadstore1.vhdl:349:31  */
  assign n19565_o = ~n19564_o;
  /* loadstore1.vhdl:353:52  */
  assign n19566_o = r3[283:278];
  /* loadstore1.vhdl:353:33  */
  assign n19567_o = {5'b0, n19566_o};  //  uext
  /* loadstore1.vhdl:353:31  */
  assign n19569_o = 11'b01110000000 - n19567_o;
  /* loadstore1.vhdl:354:51  */
  assign n19570_o = r3[282:278];
  /* loadstore1.vhdl:354:65  */
  assign n19572_o = n19570_o + 5'b00001;
  /* loadstore1.vhdl:349:13  */
  assign n19574_o = n19565_o ? 11'b00000000000 : n19569_o;
  /* loadstore1.vhdl:349:13  */
  assign n19576_o = n19565_o ? 5'b00000 : n19572_o;
  /* loadstore1.vhdl:347:13  */
  assign n19577_o = n19558_o ? n19563_o : n19574_o;
  /* loadstore1.vhdl:347:13  */
  assign n19579_o = n19558_o ? 5'b00000 : n19576_o;
  /* loadstore1.vhdl:345:13  */
  assign n19581_o = n19560_o ? 11'b11111111111 : n19577_o;
  /* loadstore1.vhdl:345:13  */
  assign n19583_o = n19560_o ? 5'b00000 : n19579_o;
  /* loadstore1.vhdl:356:46  */
  assign n19585_o = r3[276];
  /* loadstore1.vhdl:245:19  */
  assign n19593_o = n19583_o[1:0];
  /* loadstore1.vhdl:246:13  */
  assign n19595_o = n19593_o == 2'b00;
  /* loadstore1.vhdl:249:28  */
  assign n19596_o = n19555_o[21:0];
  /* loadstore1.vhdl:249:42  */
  assign n19598_o = {n19596_o, 1'b0};
  /* loadstore1.vhdl:248:13  */
  assign n19600_o = n19593_o == 2'b01;
  /* loadstore1.vhdl:251:28  */
  assign n19601_o = n19555_o[20:0];
  /* loadstore1.vhdl:251:42  */
  assign n19603_o = {n19601_o, 2'b00};
  /* loadstore1.vhdl:250:13  */
  assign n19605_o = n19593_o == 2'b10;
  /* loadstore1.vhdl:253:28  */
  assign n19606_o = n19555_o[19:0];
  /* loadstore1.vhdl:253:42  */
  assign n19608_o = {n19606_o, 3'b000};
  assign n19609_o = {n19605_o, n19600_o, n19595_o};
  /* loadstore1.vhdl:245:9  */
  always @*
    case (n19609_o)
      3'b100: n19610_o = n19603_o;
      3'b010: n19610_o = n19598_o;
      3'b001: n19610_o = n19555_o;
      default: n19610_o = n19608_o;
    endcase
  /* loadstore1.vhdl:255:19  */
  assign n19612_o = n19583_o[4:2];
  /* loadstore1.vhdl:256:13  */
  assign n19614_o = n19612_o == 3'b000;
  /* loadstore1.vhdl:259:27  */
  assign n19615_o = n19610_o[18:0];
  /* loadstore1.vhdl:259:41  */
  assign n19617_o = {n19615_o, 4'b0000};
  /* loadstore1.vhdl:258:13  */
  assign n19619_o = n19612_o == 3'b001;
  /* loadstore1.vhdl:261:27  */
  assign n19620_o = n19610_o[14:0];
  /* loadstore1.vhdl:261:41  */
  assign n19622_o = {n19620_o, 8'b00000000};
  /* loadstore1.vhdl:260:13  */
  assign n19624_o = n19612_o == 3'b010;
  /* loadstore1.vhdl:263:27  */
  assign n19625_o = n19610_o[10:0];
  /* loadstore1.vhdl:263:41  */
  assign n19627_o = {n19625_o, 12'b000000000000};
  /* loadstore1.vhdl:262:13  */
  assign n19629_o = n19612_o == 3'b011;
  /* loadstore1.vhdl:265:27  */
  assign n19630_o = n19610_o[6:0];
  /* loadstore1.vhdl:265:40  */
  assign n19632_o = {n19630_o, 16'b0000000000000000};
  /* loadstore1.vhdl:264:13  */
  assign n19634_o = n19612_o == 3'b100;
  /* loadstore1.vhdl:267:27  */
  assign n19635_o = n19610_o[2:0];
  /* loadstore1.vhdl:267:40  */
  assign n19637_o = {n19635_o, 20'b00000000000000000000};
  assign n19638_o = {n19634_o, n19629_o, n19624_o, n19619_o, n19614_o};
  /* loadstore1.vhdl:255:9  */
  always @*
    case (n19638_o)
      5'b10000: n19639_o = n19632_o;
      5'b01000: n19639_o = n19627_o;
      5'b00100: n19639_o = n19622_o;
      5'b00010: n19639_o = n19617_o;
      5'b00001: n19639_o = n19610_o;
      default: n19639_o = n19637_o;
    endcase
  /* loadstore1.vhdl:377:67  */
  assign n19654_o = n19326_o[102:71];
  /* common.vhdl:708:40  */
  assign n19659_o = n19654_o[15:11];
  /* common.vhdl:708:61  */
  assign n19660_o = n19654_o[20:16];
  /* common.vhdl:708:55  */
  assign n19661_o = {n19659_o, n19660_o};
  /* loadstore1.vhdl:379:25  */
  assign n19664_o = n19326_o[0];
  /* loadstore1.vhdl:380:29  */
  assign n19667_o = n19326_o[105:103];
  /* loadstore1.vhdl:381:30  */
  assign n19670_o = n19326_o[322];
  assign n19672_o = n19665_o[12:1];
  /* loadstore1.vhdl:382:29  */
  assign n19673_o = n19326_o[304:298];
  /* loadstore1.vhdl:383:26  */
  assign n19675_o = n19326_o[308:305];
  /* loadstore1.vhdl:384:30  */
  assign n19677_o = n19326_o[308:305];
  /* loadstore1.vhdl:385:32  */
  assign n19679_o = n19326_o[310];
  /* loadstore1.vhdl:386:31  */
  assign n19681_o = n19326_o[311];
  assign n19683_o = n19665_o[179:177];
  /* loadstore1.vhdl:387:26  */
  assign n19684_o = n19326_o[312];
  /* loadstore1.vhdl:388:24  */
  assign n19686_o = n19326_o[317:313];
  /* loadstore1.vhdl:389:27  */
  assign n19688_o = n19326_o[318];
  /* loadstore1.vhdl:390:22  */
  assign n19690_o = n19326_o[319];
  assign n19692_o = n19665_o[189:188];
  /* loadstore1.vhdl:391:22  */
  assign n19693_o = n19326_o[309];
  /* loadstore1.vhdl:392:29  */
  assign n19695_o = n19326_o[320];
  /* loadstore1.vhdl:393:29  */
  assign n19697_o = n19326_o[321];
  /* fpu.vhdl:489:18  */
  assign n19700_o = n19665_o[194];
  /* loadstore1.vhdl:395:23  */
  assign n19701_o = n19326_o[70:7];
  /* fpu.vhdl:488:18  */
  assign n19702_o = n19665_o[208:205];
  /* loadstore1.vhdl:397:52  */
  assign n19703_o = n19326_o[169:106];
  /* loadstore1.vhdl:397:75  */
  assign n19704_o = n19326_o[233:170];
  /* loadstore1.vhdl:397:59  */
  assign n19705_o = n19703_o + n19704_o;
  /* loadstore1.vhdl:399:29  */
  assign n19706_o = n19326_o[323];
  /* loadstore1.vhdl:399:20  */
  assign n19708_o = 1'b1 & n19706_o;
  /* loadstore1.vhdl:400:41  */
  assign n19710_o = {32'b00000000000000000000000000000000, store_sp_data};
  /* loadstore1.vhdl:402:34  */
  assign n19711_o = n19326_o[297:234];
  /* loadstore1.vhdl:399:9  */
  assign n19712_o = n19708_o ? n19710_o : n19711_o;
  /* loadstore1.vhdl:406:17  */
  assign n19714_o = n19326_o[325];
  /* loadstore1.vhdl:407:21  */
  assign n19715_o = n19326_o[312];
  /* loadstore1.vhdl:407:28  */
  assign n19716_o = ~n19715_o;
  /* loadstore1.vhdl:410:60  */
  assign n19717_o = r1[337:277];
  /* loadstore1.vhdl:410:75  */
  assign n19719_o = n19717_o + 61'b0000000000000000000000000000000000000000000000000000000000001;
  /* loadstore1.vhdl:410:90  */
  assign n19720_o = r1[276:274];
  /* loadstore1.vhdl:410:80  */
  assign n19721_o = {n19719_o, n19720_o};
  /* loadstore1.vhdl:417:17  */
  assign n19725_o = n19326_o[322];
  assign n19727_o = n19721_o[63:32];
  /* insn_helpers.vhdl:45:14  */
  assign n19728_o = r1[337:306];
  /* loadstore1.vhdl:407:13  */
  assign n19729_o = n19716_o ? n19727_o : n19728_o;
  assign n19730_o = n19705_o[63:32];
  /* loadstore1.vhdl:406:9  */
  assign n19731_o = n19714_o ? n19729_o : n19730_o;
  /* loadstore1.vhdl:417:9  */
  assign n19732_o = n19725_o ? 32'b00000000000000000000000000000000 : n19731_o;
  assign n19733_o = n19721_o[31:0];
  /* insn_helpers.vhdl:45:14  */
  assign n19734_o = r1[305:274];
  /* loadstore1.vhdl:407:13  */
  assign n19735_o = n19716_o ? n19733_o : n19734_o;
  assign n19736_o = n19705_o[31:0];
  /* loadstore1.vhdl:406:9  */
  assign n19737_o = n19714_o ? n19735_o : n19736_o;
  /* fpu.vhdl:999:25  */
  assign n19738_o = {n19732_o, n19737_o};
  assign n19739_o = n19665_o[93:78];
  /* insn_helpers.vhdl:45:14  */
  assign n19740_o = {n19732_o, n19737_o};
  /* loadstore1.vhdl:424:16  */
  assign n19741_o = n19740_o[31:28];
  /* loadstore1.vhdl:424:31  */
  assign n19743_o = n19741_o == 4'b1100;
  /* loadstore1.vhdl:424:49  */
  assign n19744_o = n19326_o[320];
  /* loadstore1.vhdl:424:59  */
  assign n19745_o = ~n19744_o;
  /* loadstore1.vhdl:424:40  */
  assign n19746_o = n19743_o & n19745_o;
  /* loadstore1.vhdl:424:9  */
  assign n19748_o = n19746_o ? 1'b1 : n19693_o;
  /* loadstore1.vhdl:428:60  */
  assign n19749_o = n19326_o[307:305];
  /* loadstore1.vhdl:428:74  */
  assign n19751_o = n19749_o - 3'b001;
  /* insn_helpers.vhdl:45:14  */
  assign n19753_o = {n19701_o, n19702_o, n19661_o, n19700_o, n19697_o, n19695_o, n19748_o, n19690_o, n19692_o, n19688_o, n19686_o, n19684_o, n19681_o, n19683_o, n19679_o, n19677_o, n19675_o, n19673_o, n19667_o, n19712_o, n19739_o, n19738_o, n19670_o, n19672_o, n19664_o};
  /* loadstore1.vhdl:431:37  */
  assign n19754_o = n19753_o[171:168];
  assign n19755_o = {n19732_o, n19737_o};
  /* loadstore1.vhdl:431:49  */
  assign n19756_o = n19755_o[2:0];
  /* loadstore1.vhdl:180:13  */
  assign n19769_o = n19754_o == 4'b0001;
  /* loadstore1.vhdl:182:13  */
  assign n19772_o = n19754_o == 4'b0010;
  /* loadstore1.vhdl:184:13  */
  assign n19775_o = n19754_o == 4'b0100;
  /* loadstore1.vhdl:186:13  */
  assign n19778_o = n19754_o == 4'b1000;
  /* fpu.vhdl:885:21  */
  assign n19780_o = {n19778_o, n19775_o, n19772_o, n19769_o};
  /* loadstore1.vhdl:179:9  */
  always @*
    case (n19780_o)
      4'b1000: n19781_o = 8'b11111111;
      4'b0100: n19781_o = 8'b00001111;
      4'b0010: n19781_o = 8'b00000011;
      4'b0001: n19781_o = 8'b00000001;
      default: n19781_o = 8'b00000000;
    endcase
  /* loadstore1.vhdl:201:31  */
  assign n19783_o = {8'b00000000, n19781_o};
  /* loadstore1.vhdl:203:45  */
  assign n19785_o = {28'b0, n19756_o};  //  uext
  /* loadstore1.vhdl:202:34  */
  assign n19786_o = n19783_o << n19785_o;
  /* loadstore1.vhdl:432:31  */
  assign n19787_o = n19786_o[7:0];
  /* loadstore1.vhdl:433:35  */
  assign n19789_o = n19786_o[15:8];
  /* loadstore1.vhdl:434:20  */
  assign n19790_o = n19786_o[15:8];
  /* loadstore1.vhdl:434:34  */
  assign n19792_o = n19790_o != 8'b00000000;
  assign n19794_o = n19665_o[208];
  /* loadstore1.vhdl:434:9  */
  assign n19795_o = n19792_o ? 1'b1 : n19794_o;
  assign n19797_o = {n19732_o, n19737_o};
  /* loadstore1.vhdl:439:45  */
  assign n19798_o = n19797_o[2:0];
  /* loadstore1.vhdl:439:37  */
  assign n19799_o = n19751_o & n19798_o;
  /* loadstore1.vhdl:439:23  */
  assign n19800_o = |(n19799_o);
  /* loadstore1.vhdl:440:30  */
  assign n19801_o = n19326_o[318];
  /* loadstore1.vhdl:440:38  */
  assign n19802_o = n19801_o & n19800_o;
  assign n19803_o = n19665_o[207];
  assign n19804_o = n19665_o[205];
  /* loadstore1.vhdl:441:17  */
  assign n19805_o = n19326_o[324];
  /* loadstore1.vhdl:441:39  */
  assign n19806_o = n19326_o[325];
  /* loadstore1.vhdl:441:46  */
  assign n19807_o = ~n19806_o;
  /* loadstore1.vhdl:441:30  */
  assign n19808_o = n19805_o & n19807_o;
  /* loadstore1.vhdl:441:61  */
  assign n19809_o = n19326_o[312];
  /* loadstore1.vhdl:441:68  */
  assign n19810_o = ~n19809_o;
  /* loadstore1.vhdl:441:52  */
  assign n19811_o = n19808_o & n19810_o;
  assign n19812_o = {n19732_o, n19737_o};
  /* loadstore1.vhdl:441:82  */
  assign n19813_o = n19812_o[3];
  /* loadstore1.vhdl:441:74  */
  assign n19814_o = n19811_o & n19813_o;
  /* loadstore1.vhdl:448:21  */
  assign n19815_o = n19326_o[318];
  /* loadstore1.vhdl:448:44  */
  assign n19816_o = n19326_o[6:1];
  /* loadstore1.vhdl:448:47  */
  assign n19818_o = n19816_o == 6'b011111;
  /* loadstore1.vhdl:448:66  */
  assign n19819_o = n19326_o[310];
  /* loadstore1.vhdl:448:79  */
  assign n19820_o = ~n19819_o;
  /* loadstore1.vhdl:448:57  */
  assign n19821_o = n19818_o & n19820_o;
  /* loadstore1.vhdl:448:35  */
  assign n19822_o = n19815_o | n19821_o;
  /* loadstore1.vhdl:441:9  */
  assign n19824_o = n19825_o ? 1'b1 : n19802_o;
  /* loadstore1.vhdl:441:9  */
  assign n19825_o = n19814_o & n19822_o;
  /* loadstore1.vhdl:441:9  */
  assign n19827_o = n19814_o ? 1'b1 : n19800_o;
  /* loadstore1.vhdl:453:21  */
  assign n19828_o = ~n19827_o;
  /* loadstore1.vhdl:454:26  */
  assign n19830_o = ~n19827_o;
  /* loadstore1.vhdl:454:51  */
  assign n19831_o = n19326_o[325];
  /* loadstore1.vhdl:454:70  */
  assign n19832_o = n19326_o[324];
  /* loadstore1.vhdl:454:61  */
  assign n19833_o = ~n19832_o;
  /* loadstore1.vhdl:454:58  */
  assign n19834_o = n19831_o | n19833_o;
  /* loadstore1.vhdl:454:41  */
  assign n19835_o = n19830_o & n19834_o;
  /* loadstore1.vhdl:456:19  */
  assign n19836_o = n19326_o[6:1];
  /* loadstore1.vhdl:457:13  */
  assign n19839_o = n19836_o == 6'b100000;
  /* loadstore1.vhdl:460:25  */
  assign n19840_o = n19326_o[312];
  /* loadstore1.vhdl:460:32  */
  assign n19841_o = ~n19840_o;
  /* loadstore1.vhdl:460:46  */
  assign n19842_o = n19326_o[325];
  /* loadstore1.vhdl:460:53  */
  assign n19843_o = ~n19842_o;
  /* loadstore1.vhdl:460:38  */
  assign n19844_o = n19841_o | n19843_o;
  /* loadstore1.vhdl:462:41  */
  assign n19846_o = n19326_o[323];
  /* loadstore1.vhdl:462:32  */
  assign n19848_o = 1'b1 & n19846_o;
  /* loadstore1.vhdl:460:17  */
  assign n19850_o = n19856_o ? 1'b1 : n19700_o;
  /* fpu.vhdl:412:18  */
  assign n19852_o = n19665_o[2];
  /* loadstore1.vhdl:460:17  */
  assign n19853_o = n19844_o ? 1'b1 : n19852_o;
  /* fpu.vhdl:411:18  */
  assign n19854_o = n19665_o[11];
  /* loadstore1.vhdl:460:17  */
  assign n19855_o = n19844_o ? n19854_o : 1'b1;
  /* loadstore1.vhdl:460:17  */
  assign n19856_o = n19844_o & n19848_o;
  /* loadstore1.vhdl:459:13  */
  assign n19858_o = n19836_o == 6'b011111;
  assign n19860_o = n19665_o[4:1];
  /* fpu.vhdl:421:9  */
  assign n19861_o = n19665_o[12:6];
  assign n19862_o = {n19701_o, n19795_o, n19803_o, n19824_o, n19804_o, n19661_o, n19700_o, n19697_o, n19695_o, n19748_o, n19690_o, n19835_o, n19828_o, n19688_o, n19686_o, n19684_o, n19681_o, n19683_o, n19679_o, n19677_o, n19675_o, n19673_o, n19667_o, n19712_o, n19789_o, n19787_o, n19738_o, n19670_o, n19861_o, 1'b1, n19860_o, n19664_o};
  /* loadstore1.vhdl:472:35  */
  assign n19863_o = n19862_o[191];
  /* loadstore1.vhdl:470:13  */
  assign n19865_o = n19836_o == 6'b010100;
  /* loadstore1.vhdl:475:32  */
  assign n19867_o = n19326_o[233:170];
  /* loadstore1.vhdl:476:40  */
  assign n19868_o = n19326_o[78];
  /* loadstore1.vhdl:473:13  */
  assign n19871_o = n19836_o == 6'b111000;
  /* loadstore1.vhdl:478:13  */
  assign n19874_o = n19836_o == 6'b100100;
  /* loadstore1.vhdl:482:33  */
  assign n19876_o = n19661_o[8];
  /* loadstore1.vhdl:482:44  */
  assign n19877_o = n19661_o[5];
  /* loadstore1.vhdl:482:37  */
  assign n19878_o = n19876_o | n19877_o;
  /* loadstore1.vhdl:480:13  */
  assign n19880_o = n19836_o == 6'b101000;
  /* loadstore1.vhdl:486:32  */
  assign n19882_o = n19326_o[70:7];
  /* loadstore1.vhdl:483:13  */
  assign n19885_o = n19836_o == 6'b111101;
  assign n19886_o = {n19885_o, n19880_o, n19874_o, n19871_o, n19865_o, n19858_o, n19839_o};
  /* crhelpers.vhdl:12:14  */
  assign n19887_o = n19665_o[2];
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19888_o = n19887_o;
      7'b0100000: n19888_o = n19887_o;
      7'b0010000: n19888_o = n19887_o;
      7'b0001000: n19888_o = n19887_o;
      7'b0000100: n19888_o = n19887_o;
      7'b0000010: n19888_o = n19853_o;
      7'b0000001: n19888_o = n19887_o;
      default: n19888_o = n19887_o;
    endcase
  /* insn_helpers.vhdl:22:14  */
  assign n19889_o = n19665_o[3];
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19890_o = n19889_o;
      7'b0100000: n19890_o = n19889_o;
      7'b0010000: n19890_o = n19889_o;
      7'b0001000: n19890_o = n19889_o;
      7'b0000100: n19890_o = n19889_o;
      7'b0000010: n19890_o = n19889_o;
      7'b0000001: n19890_o = 1'b1;
      default: n19890_o = n19889_o;
    endcase
  assign n19891_o = n19665_o[4];
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19892_o = n19891_o;
      7'b0100000: n19892_o = n19891_o;
      7'b0010000: n19892_o = n19891_o;
      7'b0001000: n19892_o = 1'b1;
      7'b0000100: n19892_o = n19891_o;
      7'b0000010: n19892_o = n19891_o;
      7'b0000001: n19892_o = n19891_o;
      default: n19892_o = n19891_o;
    endcase
  assign n19893_o = n19665_o[5];
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19894_o = n19893_o;
      7'b0100000: n19894_o = n19893_o;
      7'b0010000: n19894_o = n19893_o;
      7'b0001000: n19894_o = n19893_o;
      7'b0000100: n19894_o = 1'b1;
      7'b0000010: n19894_o = n19893_o;
      7'b0000001: n19894_o = n19893_o;
      default: n19894_o = n19893_o;
    endcase
  /* fpu.vhdl:642:18  */
  assign n19895_o = n19665_o[6];
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19896_o = n19895_o;
      7'b0100000: n19896_o = n19895_o;
      7'b0010000: n19896_o = 1'b1;
      7'b0001000: n19896_o = n19895_o;
      7'b0000100: n19896_o = n19895_o;
      7'b0000010: n19896_o = n19895_o;
      7'b0000001: n19896_o = n19895_o;
      default: n19896_o = n19895_o;
    endcase
  /* fpu.vhdl:641:18  */
  assign n19897_o = n19665_o[7];
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19898_o = n19897_o;
      7'b0100000: n19898_o = 1'b1;
      7'b0010000: n19898_o = n19897_o;
      7'b0001000: n19898_o = n19897_o;
      7'b0000100: n19898_o = n19897_o;
      7'b0000010: n19898_o = n19897_o;
      7'b0000001: n19898_o = n19897_o;
      default: n19898_o = n19897_o;
    endcase
  /* fpu.vhdl:640:18  */
  assign n19899_o = n19665_o[8];
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19900_o = 1'b1;
      7'b0100000: n19900_o = n19878_o;
      7'b0010000: n19900_o = n19899_o;
      7'b0001000: n19900_o = 1'b1;
      7'b0000100: n19900_o = n19899_o;
      7'b0000010: n19900_o = n19899_o;
      7'b0000001: n19900_o = n19899_o;
      default: n19900_o = n19899_o;
    endcase
  /* fpu.vhdl:639:18  */
  assign n19901_o = n19665_o[9];
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19902_o = 1'b1;
      7'b0100000: n19902_o = n19901_o;
      7'b0010000: n19902_o = n19901_o;
      7'b0001000: n19902_o = n19901_o;
      7'b0000100: n19902_o = n19901_o;
      7'b0000010: n19902_o = n19901_o;
      7'b0000001: n19902_o = n19901_o;
      default: n19902_o = n19901_o;
    endcase
  /* fpu.vhdl:638:18  */
  assign n19903_o = n19665_o[11];
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19904_o = n19903_o;
      7'b0100000: n19904_o = n19903_o;
      7'b0010000: n19904_o = n19903_o;
      7'b0001000: n19904_o = n19903_o;
      7'b0000100: n19904_o = n19903_o;
      7'b0000010: n19904_o = n19855_o;
      7'b0000001: n19904_o = n19903_o;
      default: n19904_o = n19903_o;
    endcase
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19905_o = n19882_o;
      7'b0100000: n19905_o = n19738_o;
      7'b0010000: n19905_o = n19738_o;
      7'b0001000: n19905_o = n19867_o;
      7'b0000100: n19905_o = n19738_o;
      7'b0000010: n19905_o = n19738_o;
      7'b0000001: n19905_o = n19738_o;
      default: n19905_o = n19738_o;
    endcase
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19906_o = n19700_o;
      7'b0100000: n19906_o = n19700_o;
      7'b0010000: n19906_o = n19700_o;
      7'b0001000: n19906_o = n19700_o;
      7'b0000100: n19906_o = n19700_o;
      7'b0000010: n19906_o = n19850_o;
      7'b0000001: n19906_o = n19700_o;
      default: n19906_o = n19700_o;
    endcase
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19907_o = n19804_o;
      7'b0100000: n19907_o = n19804_o;
      7'b0010000: n19907_o = n19804_o;
      7'b0001000: n19907_o = n19868_o;
      7'b0000100: n19907_o = n19804_o;
      7'b0000010: n19907_o = n19804_o;
      7'b0000001: n19907_o = n19804_o;
      default: n19907_o = n19804_o;
    endcase
  /* loadstore1.vhdl:456:9  */
  always @*
    case (n19886_o)
      7'b1000000: n19908_o = n19824_o;
      7'b0100000: n19908_o = n19824_o;
      7'b0010000: n19908_o = n19824_o;
      7'b0001000: n19908_o = n19824_o;
      7'b0000100: n19908_o = n19863_o;
      7'b0000010: n19908_o = n19824_o;
      7'b0000001: n19908_o = n19824_o;
      default: n19908_o = n19824_o;
    endcase
  assign n19910_o = n19665_o[1];
  assign n19918_o = n19665_o[12];
  /* fpu.vhdl:630:18  */
  assign n19919_o = n19665_o[10];
  /* loadstore1.vhdl:490:26  */
  assign n19920_o = n19326_o[0];
  /* fpu.vhdl:629:18  */
  assign n19921_o = {n19701_o, n19795_o, n19803_o, n19908_o, n19907_o, n19661_o, n19906_o, n19697_o, n19695_o, n19748_o, n19690_o, n19835_o, n19828_o, n19688_o, n19686_o, n19684_o, n19681_o, n19683_o, n19679_o, n19677_o, n19675_o, n19673_o, n19667_o, n19712_o, n19789_o, n19787_o, n19905_o, n19670_o, n19918_o, n19904_o, n19919_o, n19902_o, n19900_o, n19898_o, n19896_o, n19894_o, n19892_o, n19890_o, n19888_o, n19910_o, n19664_o};
  /* loadstore1.vhdl:490:39  */
  assign n19922_o = n19921_o[2];
  /* fpu.vhdl:628:18  */
  assign n19923_o = {n19701_o, n19795_o, n19803_o, n19908_o, n19907_o, n19661_o, n19906_o, n19697_o, n19695_o, n19748_o, n19690_o, n19835_o, n19828_o, n19688_o, n19686_o, n19684_o, n19681_o, n19683_o, n19679_o, n19677_o, n19675_o, n19673_o, n19667_o, n19712_o, n19789_o, n19787_o, n19905_o, n19670_o, n19918_o, n19904_o, n19919_o, n19902_o, n19900_o, n19898_o, n19896_o, n19894_o, n19892_o, n19890_o, n19888_o, n19910_o, n19664_o};
  /* loadstore1.vhdl:490:49  */
  assign n19924_o = n19923_o[3];
  /* loadstore1.vhdl:490:44  */
  assign n19925_o = n19922_o | n19924_o;
  /* execute1.vhdl:150:12  */
  assign n19926_o = {n19701_o, n19795_o, n19803_o, n19908_o, n19907_o, n19661_o, n19906_o, n19697_o, n19695_o, n19748_o, n19690_o, n19835_o, n19828_o, n19688_o, n19686_o, n19684_o, n19681_o, n19683_o, n19679_o, n19677_o, n19675_o, n19673_o, n19667_o, n19712_o, n19789_o, n19787_o, n19905_o, n19670_o, n19918_o, n19904_o, n19919_o, n19902_o, n19900_o, n19898_o, n19896_o, n19894_o, n19892_o, n19890_o, n19888_o, n19910_o, n19664_o};
  /* loadstore1.vhdl:490:60  */
  assign n19927_o = n19926_o[5];
  /* loadstore1.vhdl:490:55  */
  assign n19928_o = n19925_o | n19927_o;
  /* loadstore1.vhdl:490:32  */
  assign n19929_o = n19920_o & n19928_o;
  /* execute1.vhdl:424:18  */
  assign n19930_o = {n19701_o, n19795_o, n19803_o, n19908_o, n19907_o, n19661_o, n19906_o, n19697_o, n19695_o, n19748_o, n19690_o, n19835_o, n19828_o, n19688_o, n19686_o, n19684_o, n19681_o, n19683_o, n19679_o, n19677_o, n19675_o, n19673_o, n19667_o, n19712_o, n19789_o, n19787_o, n19905_o, n19670_o, n19918_o, n19904_o, n19919_o, n19902_o, n19900_o, n19898_o, n19896_o, n19894_o, n19892_o, n19890_o, n19888_o, n19910_o, n19664_o};
  /* loadstore1.vhdl:490:76  */
  assign n19931_o = n19930_o[206];
  /* loadstore1.vhdl:490:70  */
  assign n19932_o = ~n19931_o;
  /* loadstore1.vhdl:490:66  */
  assign n19933_o = n19929_o & n19932_o;
  /* execute1.vhdl:426:18  */
  assign n19934_o = {n19701_o, n19795_o, n19803_o, n19908_o, n19907_o, n19661_o, n19906_o, n19697_o, n19695_o, n19748_o, n19690_o, n19835_o, n19828_o, n19688_o, n19686_o, n19684_o, n19681_o, n19683_o, n19679_o, n19677_o, n19675_o, n19673_o, n19667_o, n19712_o, n19789_o, n19787_o, n19905_o, n19670_o, n19918_o, n19904_o, n19919_o, n19902_o, n19900_o, n19898_o, n19896_o, n19894_o, n19892_o, n19890_o, n19888_o, n19933_o, n19664_o};
  /* loadstore1.vhdl:494:14  */
  assign n19935_o = n19934_o[176];
  /* execute1.vhdl:427:18  */
  assign n19936_o = {n19701_o, n19795_o, n19803_o, n19908_o, n19907_o, n19661_o, n19906_o, n19697_o, n19695_o, n19748_o, n19690_o, n19835_o, n19828_o, n19688_o, n19686_o, n19684_o, n19681_o, n19683_o, n19679_o, n19677_o, n19675_o, n19673_o, n19667_o, n19712_o, n19789_o, n19787_o, n19905_o, n19670_o, n19918_o, n19904_o, n19919_o, n19902_o, n19900_o, n19898_o, n19896_o, n19894_o, n19892_o, n19890_o, n19888_o, n19933_o, n19664_o};
  /* loadstore1.vhdl:495:44  */
  assign n19937_o = n19936_o[170:168];
  /* loadstore1.vhdl:495:58  */
  assign n19939_o = n19937_o - 3'b001;
  /* loadstore1.vhdl:494:9  */
  assign n19941_o = n19935_o ? n19939_o : 3'b000;
  /* fpu.vhdl:618:18  */
  assign n19943_o = {n19701_o, n19795_o, n19803_o, n19908_o, n19907_o, n19661_o, n19906_o, n19697_o, n19695_o, n19748_o, n19690_o, n19835_o, n19828_o, n19688_o, n19686_o, n19684_o, n19681_o, n19941_o, n19679_o, n19677_o, n19675_o, n19673_o, n19667_o, n19712_o, n19789_o, n19787_o, n19905_o, n19670_o, n19918_o, n19904_o, n19919_o, n19902_o, n19900_o, n19898_o, n19896_o, n19894_o, n19892_o, n19890_o, n19888_o, n19933_o, n19664_o};
  /* loadstore1.vhdl:502:16  */
  assign n19948_o = r1[272:0];
  /* loadstore1.vhdl:502:20  */
  assign n19949_o = n19948_o[0];
  /* loadstore1.vhdl:502:35  */
  assign n19950_o = r1[272:0];
  /* loadstore1.vhdl:502:39  */
  assign n19951_o = n19950_o[1];
  /* loadstore1.vhdl:502:57  */
  assign n19952_o = r1[273];
  /* loadstore1.vhdl:502:50  */
  assign n19953_o = ~n19952_o;
  /* loadstore1.vhdl:502:46  */
  assign n19954_o = n19951_o & n19953_o;
  /* loadstore1.vhdl:503:35  */
  assign n19955_o = r1[273];
  /* loadstore1.vhdl:503:51  */
  assign n19956_o = n19358_o[66];
  /* loadstore1.vhdl:503:42  */
  assign n19957_o = n19955_o & n19956_o;
  /* loadstore1.vhdl:502:65  */
  assign n19958_o = n19954_o | n19957_o;
  /* loadstore1.vhdl:503:58  */
  assign n19959_o = n19958_o | stage2_busy_next;
  /* loadstore1.vhdl:505:35  */
  assign n19960_o = r1[272:0];
  /* loadstore1.vhdl:505:39  */
  assign n19961_o = n19960_o[1];
  /* loadstore1.vhdl:505:53  */
  assign n19962_o = r1[272:0];
  /* loadstore1.vhdl:505:57  */
  assign n19963_o = n19962_o[208];
  /* loadstore1.vhdl:505:46  */
  assign n19964_o = n19961_o & n19963_o;
  /* loadstore1.vhdl:505:79  */
  assign n19965_o = r1[272:0];
  /* loadstore1.vhdl:505:83  */
  assign n19966_o = n19965_o[207];
  /* loadstore1.vhdl:505:72  */
  assign n19967_o = ~n19966_o;
  /* loadstore1.vhdl:505:68  */
  assign n19968_o = n19964_o & n19967_o;
  /* loadstore1.vhdl:504:48  */
  assign n19969_o = n19959_o | n19968_o;
  /* loadstore1.vhdl:502:26  */
  assign n19970_o = n19949_o & n19969_o;
  /* loadstore1.vhdl:506:20  */
  assign n19971_o = r2[307];
  /* loadstore1.vhdl:506:37  */
  assign n19972_o = r2[305];
  /* loadstore1.vhdl:506:54  */
  assign n19973_o = n19358_o[0];
  /* loadstore1.vhdl:506:45  */
  assign n19974_o = n19972_o & n19973_o;
  /* loadstore1.vhdl:506:30  */
  assign n19975_o = n19971_o | n19974_o;
  /* loadstore1.vhdl:507:21  */
  assign n19976_o = r2[306];
  /* loadstore1.vhdl:507:39  */
  assign n19977_o = n19370_o[0];
  /* loadstore1.vhdl:507:30  */
  assign n19978_o = n19976_o & n19977_o;
  /* loadstore1.vhdl:506:61  */
  assign n19979_o = n19975_o | n19978_o;
  /* loadstore1.vhdl:507:51  */
  assign n19980_o = r3[84];
  /* loadstore1.vhdl:507:45  */
  assign n19981_o = n19979_o | n19980_o;
  /* loadstore1.vhdl:508:23  */
  assign n19982_o = r1[272:0];
  /* loadstore1.vhdl:508:27  */
  assign n19983_o = n19982_o[0];
  /* loadstore1.vhdl:508:40  */
  assign n19984_o = r2[272:0];
  /* loadstore1.vhdl:508:44  */
  assign n19985_o = n19984_o[0];
  /* loadstore1.vhdl:508:54  */
  assign n19986_o = ~complete;
  /* loadstore1.vhdl:508:50  */
  assign n19987_o = n19985_o & n19986_o;
  /* loadstore1.vhdl:508:33  */
  assign n19988_o = n19983_o | n19987_o;
  /* loadstore1.vhdl:510:31  */
  assign n19989_o = r3[284];
  /* loadstore1.vhdl:510:53  */
  assign n19990_o = r1[272:0];
  /* loadstore1.vhdl:510:57  */
  assign n19991_o = n19990_o[0];
  /* loadstore1.vhdl:510:70  */
  assign n19992_o = r1[272:0];
  /* loadstore1.vhdl:510:74  */
  assign n19993_o = n19992_o[8];
  /* loadstore1.vhdl:510:63  */
  assign n19994_o = n19991_o & n19993_o;
  /* loadstore1.vhdl:510:45  */
  assign n19995_o = ~n19994_o;
  /* loadstore1.vhdl:510:41  */
  assign n19996_o = n19989_o & n19995_o;
  /* loadstore1.vhdl:511:36  */
  assign n19997_o = r2[272:0];
  /* loadstore1.vhdl:511:40  */
  assign n19998_o = n19997_o[0];
  /* loadstore1.vhdl:511:53  */
  assign n19999_o = r2[272:0];
  /* loadstore1.vhdl:511:57  */
  assign n20000_o = n19999_o[8];
  /* loadstore1.vhdl:511:46  */
  assign n20001_o = n19998_o & n20000_o;
  /* loadstore1.vhdl:511:28  */
  assign n20002_o = ~n20001_o;
  /* loadstore1.vhdl:510:82  */
  assign n20003_o = n19996_o & n20002_o;
  /* loadstore1.vhdl:523:17  */
  assign n20009_o = ~busy;
  assign n20012_o = req_in[1];
  /* loadstore1.vhdl:526:13  */
  assign n20013_o = flushing ? 1'b0 : n20012_o;
  assign n20014_o = req_in[272:2];
  assign n20015_o = req_in[0];
  /* loadstore1.vhdl:532:27  */
  assign n20016_o = n19326_o[0];
  assign n20017_o = {n20014_o, n20013_o, n20015_o};
  /* loadstore1.vhdl:532:41  */
  assign n20018_o = n20017_o[1];
  /* loadstore1.vhdl:532:33  */
  assign n20019_o = n20016_o & n20018_o;
  /* loadstore1.vhdl:533:21  */
  assign n20020_o = n19326_o[0];
  assign n20021_o = {n20014_o, n20013_o, n20015_o};
  /* loadstore1.vhdl:534:32  */
  assign n20022_o = n20021_o[77:14];
  assign n20023_o = r1[337:274];
  /* loadstore1.vhdl:533:13  */
  assign n20024_o = n20020_o ? n20022_o : n20023_o;
  assign n20026_o = {n20024_o, 1'b0};
  assign n20030_o = {n20014_o, n20013_o, n20015_o};
  /* loadstore1.vhdl:523:9  */
  assign n20033_o = n20009_o ? n20019_o : 1'b0;
  /* loadstore1.vhdl:540:15  */
  assign n20035_o = r1[272:0];
  /* loadstore1.vhdl:540:19  */
  assign n20036_o = n20035_o[0];
  /* loadstore1.vhdl:541:19  */
  assign n20037_o = r1[272:0];
  /* loadstore1.vhdl:541:23  */
  assign n20038_o = n20037_o[1];
  /* loadstore1.vhdl:541:43  */
  assign n20039_o = r1[273];
  /* loadstore1.vhdl:541:50  */
  assign n20040_o = ~n20039_o;
  /* loadstore1.vhdl:541:36  */
  assign n20041_o = n20038_o & n20040_o;
  /* loadstore1.vhdl:543:22  */
  assign n20042_o = r1[273];
  /* loadstore1.vhdl:543:44  */
  assign n20043_o = n19358_o[66];
  /* loadstore1.vhdl:543:35  */
  assign n20044_o = n20042_o & n20043_o;
  /* loadstore1.vhdl:545:36  */
  assign n20046_o = ~stage2_busy_next;
  /* loadstore1.vhdl:548:23  */
  assign n20047_o = r1[272:0];
  /* loadstore1.vhdl:548:27  */
  assign n20048_o = n20047_o[1];
  /* loadstore1.vhdl:548:47  */
  assign n20049_o = r1[272:0];
  /* loadstore1.vhdl:548:51  */
  assign n20050_o = n20049_o[208];
  /* loadstore1.vhdl:548:40  */
  assign n20051_o = n20048_o & n20050_o;
  /* loadstore1.vhdl:548:75  */
  assign n20052_o = r1[272:0];
  /* loadstore1.vhdl:548:79  */
  assign n20053_o = n20052_o[207];
  /* loadstore1.vhdl:548:91  */
  assign n20054_o = ~n20053_o;
  /* loadstore1.vhdl:548:68  */
  assign n20055_o = n20051_o & n20054_o;
  /* loadstore1.vhdl:551:71  */
  assign n20057_o = r1[77:17];
  /* loadstore1.vhdl:551:86  */
  assign n20059_o = n20057_o + 61'b0000000000000000000000000000000000000000000000000000000000001;
  /* loadstore1.vhdl:551:91  */
  assign n20061_o = {n20059_o, 3'b000};
  /* loadstore1.vhdl:552:27  */
  assign n20062_o = r1[272:0];
  /* loadstore1.vhdl:552:31  */
  assign n20063_o = n20062_o[13];
  assign n20065_o = n20061_o[32];
  /* loadstore1.vhdl:552:21  */
  assign n20066_o = n20063_o ? 1'b0 : n20065_o;
  assign n20067_o = n20061_o[63:33];
  assign n20068_o = n20061_o[31:0];
  /* loadstore1.vhdl:555:40  */
  assign n20069_o = r1[272:0];
  /* loadstore1.vhdl:555:44  */
  assign n20070_o = n20069_o[93:86];
  assign n20071_o = {n20070_o, n20067_o, n20066_o, n20068_o};
  assign n20072_o = n20030_o[85:14];
  assign n20073_o = r1[85:14];
  /* loadstore1.vhdl:523:9  */
  assign n20074_o = n20009_o ? n20072_o : n20073_o;
  /* loadstore1.vhdl:548:17  */
  assign n20075_o = n20055_o ? n20071_o : n20074_o;
  assign n20076_o = n20030_o[207];
  assign n20077_o = r1[207];
  /* loadstore1.vhdl:523:9  */
  assign n20078_o = n20009_o ? n20076_o : n20077_o;
  /* loadstore1.vhdl:548:17  */
  assign n20079_o = n20055_o ? 1'b1 : n20078_o;
  /* loadstore1.vhdl:545:13  */
  assign n20081_o = n20090_o ? 1'b1 : n20033_o;
  assign n20082_o = n20030_o[85:14];
  assign n20083_o = r1[85:14];
  /* loadstore1.vhdl:523:9  */
  assign n20084_o = n20009_o ? n20082_o : n20083_o;
  /* loadstore1.vhdl:545:13  */
  assign n20085_o = n20046_o ? n20075_o : n20084_o;
  assign n20086_o = n20030_o[207];
  assign n20087_o = r1[207];
  /* loadstore1.vhdl:523:9  */
  assign n20088_o = n20009_o ? n20086_o : n20087_o;
  /* loadstore1.vhdl:545:13  */
  assign n20089_o = n20046_o ? n20079_o : n20088_o;
  /* loadstore1.vhdl:545:13  */
  assign n20090_o = n20046_o & n20055_o;
  assign n20091_o = n20026_o[0];
  assign n20092_o = r1[273];
  /* loadstore1.vhdl:523:9  */
  assign n20093_o = n20009_o ? n20091_o : n20092_o;
  /* loadstore1.vhdl:543:13  */
  assign n20094_o = n20044_o ? 1'b0 : n20093_o;
  assign n20095_o = n20030_o[85:14];
  assign n20096_o = r1[85:14];
  /* loadstore1.vhdl:523:9  */
  assign n20097_o = n20009_o ? n20095_o : n20096_o;
  /* loadstore1.vhdl:543:13  */
  assign n20098_o = n20044_o ? n20097_o : n20085_o;
  assign n20099_o = n20030_o[207];
  assign n20100_o = r1[207];
  /* loadstore1.vhdl:523:9  */
  assign n20101_o = n20009_o ? n20099_o : n20100_o;
  /* loadstore1.vhdl:543:13  */
  assign n20102_o = n20044_o ? n20101_o : n20089_o;
  /* loadstore1.vhdl:543:13  */
  assign n20103_o = n20044_o ? n20033_o : n20081_o;
  assign n20104_o = n20026_o[0];
  assign n20105_o = r1[273];
  /* loadstore1.vhdl:523:9  */
  assign n20106_o = n20009_o ? n20104_o : n20105_o;
  /* loadstore1.vhdl:541:13  */
  assign n20107_o = n20041_o ? n20106_o : n20094_o;
  assign n20108_o = n20030_o[85:14];
  assign n20109_o = r1[85:14];
  /* loadstore1.vhdl:523:9  */
  assign n20110_o = n20009_o ? n20108_o : n20109_o;
  /* loadstore1.vhdl:541:13  */
  assign n20111_o = n20041_o ? n20110_o : n20098_o;
  assign n20112_o = n20030_o[207];
  assign n20113_o = r1[207];
  /* loadstore1.vhdl:523:9  */
  assign n20114_o = n20009_o ? n20112_o : n20113_o;
  /* loadstore1.vhdl:541:13  */
  assign n20115_o = n20041_o ? n20114_o : n20102_o;
  /* loadstore1.vhdl:541:13  */
  assign n20117_o = n20041_o ? 1'b1 : n20103_o;
  assign n20118_o = n20026_o[0];
  assign n20119_o = r1[273];
  /* loadstore1.vhdl:523:9  */
  assign n20120_o = n20009_o ? n20118_o : n20119_o;
  /* loadstore1.vhdl:540:9  */
  assign n20121_o = n20036_o ? n20107_o : n20120_o;
  assign n20122_o = n20026_o[64:1];
  assign n20123_o = r1[337:274];
  /* loadstore1.vhdl:523:9  */
  assign n20124_o = n20009_o ? n20122_o : n20123_o;
  assign n20125_o = n20030_o[85:14];
  assign n20126_o = r1[85:14];
  /* loadstore1.vhdl:523:9  */
  assign n20127_o = n20009_o ? n20125_o : n20126_o;
  /* loadstore1.vhdl:540:9  */
  assign n20128_o = n20036_o ? n20111_o : n20127_o;
  assign n20129_o = n20030_o[207];
  assign n20130_o = r1[207];
  /* loadstore1.vhdl:523:9  */
  assign n20131_o = n20009_o ? n20129_o : n20130_o;
  /* loadstore1.vhdl:540:9  */
  assign n20132_o = n20036_o ? n20115_o : n20131_o;
  assign n20139_o = n20030_o[272:208];
  assign n20140_o = r1[272:208];
  /* loadstore1.vhdl:523:9  */
  assign n20141_o = n20009_o ? n20139_o : n20140_o;
  assign n20142_o = n20030_o[206:86];
  assign n20143_o = r1[206:86];
  /* loadstore1.vhdl:523:9  */
  assign n20144_o = n20009_o ? n20142_o : n20143_o;
  /* loadstore1.vhdl:540:9  */
  assign n20145_o = n20036_o ? n20117_o : n20033_o;
  /* loadstore1.vhdl:560:17  */
  assign n20146_o = r3in[285];
  assign n20148_o = n20030_o[0];
  assign n20149_o = r1[0];
  /* loadstore1.vhdl:523:9  */
  assign n20150_o = n20009_o ? n20148_o : n20149_o;
  /* loadstore1.vhdl:560:9  */
  assign n20151_o = n20146_o ? 1'b0 : n20150_o;
  assign n20152_o = n20030_o[13:1];
  assign n20153_o = r1[13:1];
  /* loadstore1.vhdl:523:9  */
  assign n20154_o = n20009_o ? n20152_o : n20153_o;
  /* loadstore1.vhdl:560:9  */
  assign n20156_o = n20146_o ? 1'b0 : n20145_o;
  assign n20157_o = {n20141_o, n20132_o, n20144_o, n20128_o, n20154_o, n20151_o};
  /* loadstore1.vhdl:566:24  */
  assign n20158_o = n20156_o & stage1_issue_enable;
  /* loadstore1.vhdl:566:61  */
  assign n20159_o = n19358_o[66];
  /* loadstore1.vhdl:566:52  */
  assign n20160_o = ~n20159_o;
  /* loadstore1.vhdl:566:48  */
  assign n20161_o = n20158_o & n20160_o;
  /* loadstore1.vhdl:566:71  */
  assign n20162_o = ~dc_stall;
  /* loadstore1.vhdl:566:67  */
  assign n20163_o = n20161_o & n20162_o;
  /* loadstore1.vhdl:567:9  */
  assign n20164_o = n20156_o ? n20163_o : n20121_o;
  assign n20165_o = {n20141_o, n20132_o, n20144_o, n20128_o, n20154_o, n20151_o};
  assign n20166_o = {n20124_o, n20164_o, n20157_o};
  /* loadstore1.vhdl:591:41  */
  assign n20177_o = r1[276:274];
  /* loadstore1.vhdl:593:37  */
  assign n20179_o = 3'b000 - n20177_o;
  /* loadstore1.vhdl:593:59  */
  assign n20180_o = r1[272:0];
  /* loadstore1.vhdl:593:63  */
  assign n20181_o = n20180_o[179:177];
  /* loadstore1.vhdl:593:52  */
  assign n20182_o = n20179_o ^ n20181_o;
  /* loadstore1.vhdl:593:37  */
  assign n20192_o = 3'b001 - n20177_o;
  /* loadstore1.vhdl:593:59  */
  assign n20193_o = r1[272:0];
  /* loadstore1.vhdl:593:63  */
  assign n20194_o = n20193_o[179:177];
  /* loadstore1.vhdl:593:52  */
  assign n20195_o = n20192_o ^ n20194_o;
  /* loadstore1.vhdl:593:37  */
  assign n20205_o = 3'b010 - n20177_o;
  /* loadstore1.vhdl:593:59  */
  assign n20206_o = r1[272:0];
  /* loadstore1.vhdl:593:63  */
  assign n20207_o = n20206_o[179:177];
  /* loadstore1.vhdl:593:52  */
  assign n20208_o = n20205_o ^ n20207_o;
  /* loadstore1.vhdl:593:37  */
  assign n20218_o = 3'b011 - n20177_o;
  /* loadstore1.vhdl:593:59  */
  assign n20219_o = r1[272:0];
  /* loadstore1.vhdl:593:63  */
  assign n20220_o = n20219_o[179:177];
  /* loadstore1.vhdl:593:52  */
  assign n20221_o = n20218_o ^ n20220_o;
  /* loadstore1.vhdl:593:37  */
  assign n20231_o = 3'b100 - n20177_o;
  /* loadstore1.vhdl:593:59  */
  assign n20232_o = r1[272:0];
  /* loadstore1.vhdl:593:63  */
  assign n20233_o = n20232_o[179:177];
  /* loadstore1.vhdl:593:52  */
  assign n20234_o = n20231_o ^ n20233_o;
  /* loadstore1.vhdl:593:37  */
  assign n20244_o = 3'b101 - n20177_o;
  /* loadstore1.vhdl:593:59  */
  assign n20245_o = r1[272:0];
  /* loadstore1.vhdl:593:63  */
  assign n20246_o = n20245_o[179:177];
  /* loadstore1.vhdl:593:52  */
  assign n20247_o = n20244_o ^ n20246_o;
  /* loadstore1.vhdl:593:37  */
  assign n20257_o = 3'b110 - n20177_o;
  /* loadstore1.vhdl:593:59  */
  assign n20258_o = r1[272:0];
  /* loadstore1.vhdl:593:63  */
  assign n20259_o = n20258_o[179:177];
  /* loadstore1.vhdl:593:52  */
  assign n20260_o = n20257_o ^ n20259_o;
  /* loadstore1.vhdl:593:37  */
  assign n20270_o = 3'b111 - n20177_o;
  /* loadstore1.vhdl:593:59  */
  assign n20271_o = r1[272:0];
  /* loadstore1.vhdl:593:63  */
  assign n20272_o = n20271_o[179:177];
  /* loadstore1.vhdl:593:52  */
  assign n20273_o = n20270_o ^ n20272_o;
  /* loadstore1.vhdl:598:29  */
  assign n20282_o = ~stage3_busy_next;
  /* loadstore1.vhdl:599:17  */
  assign n20283_o = r1[272:0];
  /* loadstore1.vhdl:599:21  */
  assign n20284_o = n20283_o[0];
  /* loadstore1.vhdl:599:27  */
  assign n20285_o = ~n20284_o;
  /* loadstore1.vhdl:599:39  */
  assign n20286_o = r1[273];
  /* loadstore1.vhdl:599:33  */
  assign n20287_o = n20285_o | n20286_o;
  /* loadstore1.vhdl:599:58  */
  assign n20288_o = r1[272:0];
  /* loadstore1.vhdl:599:62  */
  assign n20289_o = n20288_o[1];
  /* loadstore1.vhdl:599:69  */
  assign n20290_o = ~n20289_o;
  /* loadstore1.vhdl:599:52  */
  assign n20291_o = n20287_o | n20290_o;
  /* loadstore1.vhdl:598:35  */
  assign n20292_o = n20282_o & n20291_o;
  /* loadstore1.vhdl:601:27  */
  assign n20294_o = r1[337:274];
  assign n20295_o = r1[272:158];
  assign n20296_o = r1[93:0];
  /* loadstore1.vhdl:603:29  */
  assign n20297_o = r1[272:0];
  /* loadstore1.vhdl:603:33  */
  assign n20298_o = n20297_o[0];
  /* loadstore1.vhdl:603:46  */
  assign n20299_o = r1[272:0];
  /* loadstore1.vhdl:603:50  */
  assign n20300_o = n20299_o[1];
  /* loadstore1.vhdl:603:39  */
  assign n20301_o = n20298_o & n20300_o;
  /* loadstore1.vhdl:603:68  */
  assign n20302_o = r1[272:0];
  /* loadstore1.vhdl:603:72  */
  assign n20303_o = n20302_o[194];
  /* loadstore1.vhdl:603:61  */
  assign n20304_o = ~n20303_o;
  /* loadstore1.vhdl:603:57  */
  assign n20305_o = n20301_o & n20304_o;
  /* loadstore1.vhdl:604:34  */
  assign n20306_o = r1[272:0];
  /* loadstore1.vhdl:604:38  */
  assign n20307_o = n20306_o[208];
  /* loadstore1.vhdl:604:60  */
  assign n20308_o = r1[272:0];
  /* loadstore1.vhdl:604:64  */
  assign n20309_o = n20308_o[207];
  /* loadstore1.vhdl:604:53  */
  assign n20310_o = ~n20309_o;
  /* loadstore1.vhdl:604:49  */
  assign n20311_o = n20307_o & n20310_o;
  /* loadstore1.vhdl:604:26  */
  assign n20312_o = ~n20311_o;
  /* loadstore1.vhdl:603:80  */
  assign n20313_o = n20305_o & n20312_o;
  /* loadstore1.vhdl:605:30  */
  assign n20314_o = r1[272:0];
  /* loadstore1.vhdl:605:34  */
  assign n20315_o = n20314_o[0];
  /* loadstore1.vhdl:605:47  */
  assign n20316_o = r1[272:0];
  /* loadstore1.vhdl:605:51  */
  assign n20317_o = n20316_o[8];
  /* loadstore1.vhdl:605:40  */
  assign n20318_o = n20315_o & n20317_o;
  /* loadstore1.vhdl:606:31  */
  assign n20319_o = r1[272:0];
  /* loadstore1.vhdl:606:35  */
  assign n20320_o = n20319_o[0];
  /* loadstore1.vhdl:606:49  */
  assign n20321_o = r1[272:0];
  /* loadstore1.vhdl:606:53  */
  assign n20322_o = n20321_o[12];
  /* loadstore1.vhdl:606:64  */
  assign n20323_o = r1[272:0];
  /* loadstore1.vhdl:606:68  */
  assign n20324_o = n20323_o[6];
  /* loadstore1.vhdl:606:58  */
  assign n20325_o = n20322_o | n20324_o;
  /* loadstore1.vhdl:607:50  */
  assign n20326_o = r1[272:0];
  /* loadstore1.vhdl:607:54  */
  assign n20327_o = n20326_o[7];
  /* loadstore1.vhdl:607:75  */
  assign n20328_o = r1[272:0];
  /* loadstore1.vhdl:607:79  */
  assign n20329_o = n20328_o[8];
  /* loadstore1.vhdl:607:68  */
  assign n20330_o = ~n20329_o;
  /* loadstore1.vhdl:607:64  */
  assign n20331_o = n20327_o & n20330_o;
  /* loadstore1.vhdl:606:77  */
  assign n20332_o = n20325_o | n20331_o;
  /* loadstore1.vhdl:608:49  */
  assign n20333_o = r1[272:0];
  /* loadstore1.vhdl:608:53  */
  assign n20334_o = n20333_o[10];
  /* loadstore1.vhdl:607:87  */
  assign n20335_o = n20332_o | n20334_o;
  /* loadstore1.vhdl:608:69  */
  assign n20336_o = r1[272:0];
  /* loadstore1.vhdl:608:73  */
  assign n20337_o = n20336_o[11];
  /* loadstore1.vhdl:608:63  */
  assign n20338_o = n20335_o | n20337_o;
  /* loadstore1.vhdl:606:41  */
  assign n20339_o = n20320_o & n20338_o;
  /* loadstore1.vhdl:609:19  */
  assign n20340_o = r1[272:0];
  /* loadstore1.vhdl:609:23  */
  assign n20341_o = n20340_o[6];
  /* loadstore1.vhdl:611:22  */
  assign n20343_o = r1[272:0];
  /* loadstore1.vhdl:611:26  */
  assign n20344_o = n20343_o[11];
  /* loadstore1.vhdl:611:48  */
  assign n20345_o = r1[272:0];
  /* loadstore1.vhdl:611:52  */
  assign n20346_o = n20345_o[3];
  /* loadstore1.vhdl:611:42  */
  assign n20347_o = n20344_o | n20346_o;
  /* loadstore1.vhdl:613:22  */
  assign n20349_o = r1[272:0];
  /* loadstore1.vhdl:613:26  */
  assign n20350_o = n20349_o[194];
  /* loadstore1.vhdl:613:13  */
  assign n20353_o = n20350_o ? 2'b10 : 2'b11;
  /* loadstore1.vhdl:611:13  */
  assign n20354_o = n20347_o ? 2'b01 : n20353_o;
  /* loadstore1.vhdl:609:13  */
  assign n20355_o = n20341_o ? 2'b00 : n20354_o;
  /* loadstore1.vhdl:621:49  */
  assign n20356_o = r1[272:0];
  /* loadstore1.vhdl:621:53  */
  assign n20357_o = n20356_o[179:177];
  /* loadstore1.vhdl:621:42  */
  assign n20359_o = 3'b000 ^ n20357_o;
  /* loadstore1.vhdl:622:28  */
  assign n20361_o = {1'b0, n20359_o};
  /* loadstore1.vhdl:622:42  */
  assign n20363_o = {1'b0, n20177_o};
  /* loadstore1.vhdl:622:35  */
  assign n20364_o = n20361_o + n20363_o;
  /* loadstore1.vhdl:623:38  */
  assign n20365_o = n20364_o[3];
  /* loadstore1.vhdl:624:38  */
  assign n20366_o = n20364_o[2:0];
  /* loadstore1.vhdl:621:49  */
  assign n20367_o = r1[272:0];
  /* loadstore1.vhdl:621:53  */
  assign n20368_o = n20367_o[179:177];
  /* loadstore1.vhdl:621:42  */
  assign n20370_o = 3'b001 ^ n20368_o;
  /* loadstore1.vhdl:622:28  */
  assign n20372_o = {1'b0, n20370_o};
  /* loadstore1.vhdl:622:42  */
  assign n20374_o = {1'b0, n20177_o};
  /* loadstore1.vhdl:622:35  */
  assign n20375_o = n20372_o + n20374_o;
  /* loadstore1.vhdl:623:38  */
  assign n20376_o = n20375_o[3];
  /* loadstore1.vhdl:624:38  */
  assign n20377_o = n20375_o[2:0];
  /* loadstore1.vhdl:621:49  */
  assign n20378_o = r1[272:0];
  /* loadstore1.vhdl:621:53  */
  assign n20379_o = n20378_o[179:177];
  /* loadstore1.vhdl:621:42  */
  assign n20381_o = 3'b010 ^ n20379_o;
  /* loadstore1.vhdl:622:28  */
  assign n20383_o = {1'b0, n20381_o};
  /* loadstore1.vhdl:622:42  */
  assign n20385_o = {1'b0, n20177_o};
  /* loadstore1.vhdl:622:35  */
  assign n20386_o = n20383_o + n20385_o;
  /* loadstore1.vhdl:623:38  */
  assign n20387_o = n20386_o[3];
  /* loadstore1.vhdl:624:38  */
  assign n20388_o = n20386_o[2:0];
  /* loadstore1.vhdl:621:49  */
  assign n20389_o = r1[272:0];
  /* loadstore1.vhdl:621:53  */
  assign n20390_o = n20389_o[179:177];
  /* loadstore1.vhdl:621:42  */
  assign n20392_o = 3'b011 ^ n20390_o;
  /* loadstore1.vhdl:622:28  */
  assign n20394_o = {1'b0, n20392_o};
  /* loadstore1.vhdl:622:42  */
  assign n20396_o = {1'b0, n20177_o};
  /* loadstore1.vhdl:622:35  */
  assign n20397_o = n20394_o + n20396_o;
  /* loadstore1.vhdl:623:38  */
  assign n20398_o = n20397_o[3];
  /* loadstore1.vhdl:624:38  */
  assign n20399_o = n20397_o[2:0];
  /* loadstore1.vhdl:621:49  */
  assign n20400_o = r1[272:0];
  /* loadstore1.vhdl:621:53  */
  assign n20401_o = n20400_o[179:177];
  /* loadstore1.vhdl:621:42  */
  assign n20403_o = 3'b100 ^ n20401_o;
  /* loadstore1.vhdl:622:28  */
  assign n20405_o = {1'b0, n20403_o};
  /* loadstore1.vhdl:622:42  */
  assign n20407_o = {1'b0, n20177_o};
  /* loadstore1.vhdl:622:35  */
  assign n20408_o = n20405_o + n20407_o;
  /* loadstore1.vhdl:623:38  */
  assign n20409_o = n20408_o[3];
  /* loadstore1.vhdl:624:38  */
  assign n20410_o = n20408_o[2:0];
  /* loadstore1.vhdl:621:49  */
  assign n20411_o = r1[272:0];
  /* loadstore1.vhdl:621:53  */
  assign n20412_o = n20411_o[179:177];
  /* loadstore1.vhdl:621:42  */
  assign n20414_o = 3'b101 ^ n20412_o;
  /* loadstore1.vhdl:622:28  */
  assign n20416_o = {1'b0, n20414_o};
  /* loadstore1.vhdl:622:42  */
  assign n20418_o = {1'b0, n20177_o};
  /* loadstore1.vhdl:622:35  */
  assign n20419_o = n20416_o + n20418_o;
  /* loadstore1.vhdl:623:38  */
  assign n20420_o = n20419_o[3];
  /* loadstore1.vhdl:624:38  */
  assign n20421_o = n20419_o[2:0];
  /* loadstore1.vhdl:621:49  */
  assign n20422_o = r1[272:0];
  /* loadstore1.vhdl:621:53  */
  assign n20423_o = n20422_o[179:177];
  /* loadstore1.vhdl:621:42  */
  assign n20425_o = 3'b110 ^ n20423_o;
  /* loadstore1.vhdl:622:28  */
  assign n20427_o = {1'b0, n20425_o};
  /* loadstore1.vhdl:622:42  */
  assign n20429_o = {1'b0, n20177_o};
  /* loadstore1.vhdl:622:35  */
  assign n20430_o = n20427_o + n20429_o;
  /* loadstore1.vhdl:623:38  */
  assign n20431_o = n20430_o[3];
  /* loadstore1.vhdl:624:38  */
  assign n20432_o = n20430_o[2:0];
  /* loadstore1.vhdl:621:49  */
  assign n20433_o = r1[272:0];
  /* loadstore1.vhdl:621:53  */
  assign n20434_o = n20433_o[179:177];
  /* loadstore1.vhdl:621:42  */
  assign n20436_o = 3'b111 ^ n20434_o;
  /* loadstore1.vhdl:622:28  */
  assign n20438_o = {1'b0, n20436_o};
  /* loadstore1.vhdl:622:42  */
  assign n20440_o = {1'b0, n20177_o};
  /* loadstore1.vhdl:622:35  */
  assign n20441_o = n20438_o + n20440_o;
  /* loadstore1.vhdl:623:38  */
  assign n20442_o = n20441_o[3];
  /* loadstore1.vhdl:624:38  */
  assign n20443_o = n20441_o[2:0];
  /* loadstore1.vhdl:626:32  */
  assign n20444_o = ~stage3_busy_next;
  assign n20448_o = {1'b0, 1'b0};
  assign n20449_o = r2[0];
  /* loadstore1.vhdl:626:9  */
  assign n20450_o = n20444_o ? 1'b0 : n20449_o;
  assign n20451_o = r2[306:305];
  /* loadstore1.vhdl:626:9  */
  assign n20452_o = n20444_o ? n20448_o : n20451_o;
  assign n20453_o = {n20294_o, n20355_o, n20339_o, n20318_o, n20313_o, n20442_o, n20431_o, n20420_o, n20409_o, n20398_o, n20387_o, n20376_o, n20365_o, n20366_o, n20377_o, n20388_o, n20399_o, n20410_o, n20421_o, n20432_o, n20443_o, n20295_o, store_data, n20296_o};
  assign n20454_o = n20453_o[0];
  /* loadstore1.vhdl:598:9  */
  assign n20455_o = n20292_o ? n20454_o : n20450_o;
  assign n20456_o = n20453_o[304:1];
  assign n20457_o = r2[304:1];
  /* loadstore1.vhdl:598:9  */
  assign n20458_o = n20292_o ? n20456_o : n20457_o;
  assign n20459_o = n20453_o[306:305];
  /* loadstore1.vhdl:598:9  */
  assign n20460_o = n20292_o ? n20459_o : n20452_o;
  assign n20461_o = n20453_o[373:307];
  assign n20462_o = r2[373:307];
  /* loadstore1.vhdl:598:9  */
  assign n20463_o = n20292_o ? n20461_o : n20462_o;
  /* loadstore1.vhdl:632:32  */
  assign n20469_o = r1[272:0];
  /* loadstore1.vhdl:632:36  */
  assign n20470_o = n20469_o[0];
  /* loadstore1.vhdl:632:42  */
  assign n20471_o = n20470_o & stage3_busy_next;
  /* loadstore1.vhdl:634:17  */
  assign n20472_o = r3in[285];
  /* loadstore1.vhdl:634:9  */
  assign n20474_o = n20472_o ? 1'b0 : n20455_o;
  assign n20475_o = {n20463_o, n20460_o, n20458_o, n20474_o};
  /* loadstore1.vhdl:684:42  */
  assign n20504_o = r2[296:294];
  /* loadstore1.vhdl:684:42  */
  assign n20513_o = r2[293:291];
  /* loadstore1.vhdl:684:42  */
  assign n20522_o = r2[290:288];
  /* loadstore1.vhdl:684:42  */
  assign n20531_o = r2[287:285];
  /* loadstore1.vhdl:684:42  */
  assign n20540_o = r2[284:282];
  /* loadstore1.vhdl:684:42  */
  assign n20549_o = r2[281:279];
  /* loadstore1.vhdl:684:42  */
  assign n20558_o = r2[278:276];
  /* loadstore1.vhdl:684:42  */
  assign n20567_o = r2[275:273];
  /* loadstore1.vhdl:692:15  */
  assign n20576_o = r2[272:0];
  /* loadstore1.vhdl:692:19  */
  assign n20577_o = n20576_o[207];
  /* loadstore1.vhdl:692:44  */
  assign n20578_o = r2[272:0];
  /* loadstore1.vhdl:692:48  */
  assign n20579_o = n20578_o[176];
  /* loadstore1.vhdl:692:37  */
  assign n20580_o = n20577_o & n20579_o;
  /* loadstore1.vhdl:693:39  */
  assign n20581_o = r2[171];
  /* loadstore1.vhdl:693:59  */
  assign n20582_o = r3[148];
  /* loadstore1.vhdl:693:43  */
  assign n20583_o = n20581_o & n20582_o;
  /* loadstore1.vhdl:694:39  */
  assign n20584_o = r2[170];
  /* loadstore1.vhdl:694:59  */
  assign n20585_o = r3[116];
  /* loadstore1.vhdl:694:43  */
  assign n20586_o = n20584_o & n20585_o;
  /* loadstore1.vhdl:693:65  */
  assign n20587_o = n20583_o | n20586_o;
  /* loadstore1.vhdl:695:39  */
  assign n20588_o = r2[169];
  /* loadstore1.vhdl:695:59  */
  assign n20589_o = r3[100];
  /* loadstore1.vhdl:695:43  */
  assign n20590_o = n20588_o & n20589_o;
  /* loadstore1.vhdl:694:65  */
  assign n20591_o = n20587_o | n20590_o;
  /* loadstore1.vhdl:696:39  */
  assign n20592_o = r2[168];
  /* loadstore1.vhdl:696:59  */
  assign n20593_o = r3[92];
  /* loadstore1.vhdl:696:43  */
  assign n20594_o = n20592_o & n20593_o;
  /* loadstore1.vhdl:695:65  */
  assign n20595_o = n20591_o | n20594_o;
  /* loadstore1.vhdl:698:39  */
  assign n20596_o = r2[171];
  assign n20597_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:698:60  */
  assign n20598_o = n20597_o[63];
  /* loadstore1.vhdl:698:43  */
  assign n20599_o = n20596_o & n20598_o;
  /* loadstore1.vhdl:699:39  */
  assign n20600_o = r2[170];
  assign n20601_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:699:60  */
  assign n20602_o = n20601_o[31];
  /* loadstore1.vhdl:699:43  */
  assign n20603_o = n20600_o & n20602_o;
  /* loadstore1.vhdl:698:66  */
  assign n20604_o = n20599_o | n20603_o;
  /* loadstore1.vhdl:700:39  */
  assign n20605_o = r2[169];
  assign n20606_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:700:60  */
  assign n20607_o = n20606_o[15];
  /* loadstore1.vhdl:700:43  */
  assign n20608_o = n20605_o & n20607_o;
  /* loadstore1.vhdl:699:66  */
  assign n20609_o = n20604_o | n20608_o;
  /* loadstore1.vhdl:701:39  */
  assign n20610_o = r2[168];
  assign n20611_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:701:60  */
  assign n20612_o = n20611_o[7];
  /* loadstore1.vhdl:701:43  */
  assign n20613_o = n20610_o & n20612_o;
  /* loadstore1.vhdl:700:66  */
  assign n20614_o = n20609_o | n20613_o;
  /* loadstore1.vhdl:692:9  */
  assign n20615_o = n20580_o ? n20595_o : n20614_o;
  /* loadstore1.vhdl:706:43  */
  assign n20616_o = r2[272:0];
  /* loadstore1.vhdl:706:47  */
  assign n20617_o = n20616_o[171:168];
  /* loadstore1.vhdl:706:20  */
  assign n20618_o = {27'b0, n20617_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20619_o = {1'b0, n20618_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20621_o = $signed(32'b00000000000000000000000000000000) < $signed(n20619_o);
  /* loadstore1.vhdl:707:23  */
  assign n20622_o = r2[272:0];
  /* loadstore1.vhdl:707:27  */
  assign n20623_o = n20622_o[207];
  /* loadstore1.vhdl:708:59  */
  assign n20624_o = r2[297];
  /* loadstore1.vhdl:708:42  */
  assign n20625_o = ~n20624_o;
  /* loadstore1.vhdl:708:40  */
  assign n20627_o = {1'b1, n20625_o};
  /* loadstore1.vhdl:707:17  */
  assign n20629_o = n20623_o ? n20627_o : 2'b10;
  /* loadstore1.vhdl:706:13  */
  assign n20631_o = n20621_o ? n20629_o : 2'b00;
  /* loadstore1.vhdl:706:43  */
  assign n20632_o = r2[272:0];
  /* loadstore1.vhdl:706:47  */
  assign n20633_o = n20632_o[171:168];
  /* loadstore1.vhdl:706:20  */
  assign n20634_o = {27'b0, n20633_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20635_o = {1'b0, n20634_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20637_o = $signed(32'b00000000000000000000000000000001) < $signed(n20635_o);
  /* loadstore1.vhdl:707:23  */
  assign n20638_o = r2[272:0];
  /* loadstore1.vhdl:707:27  */
  assign n20639_o = n20638_o[207];
  /* loadstore1.vhdl:708:59  */
  assign n20640_o = r2[298];
  /* loadstore1.vhdl:708:42  */
  assign n20641_o = ~n20640_o;
  /* loadstore1.vhdl:708:40  */
  assign n20643_o = {1'b1, n20641_o};
  /* loadstore1.vhdl:707:17  */
  assign n20645_o = n20639_o ? n20643_o : 2'b10;
  /* loadstore1.vhdl:706:13  */
  assign n20647_o = n20637_o ? n20645_o : 2'b00;
  /* loadstore1.vhdl:706:43  */
  assign n20648_o = r2[272:0];
  /* loadstore1.vhdl:706:47  */
  assign n20649_o = n20648_o[171:168];
  /* loadstore1.vhdl:706:20  */
  assign n20650_o = {27'b0, n20649_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20651_o = {1'b0, n20650_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20653_o = $signed(32'b00000000000000000000000000000010) < $signed(n20651_o);
  /* loadstore1.vhdl:707:23  */
  assign n20654_o = r2[272:0];
  /* loadstore1.vhdl:707:27  */
  assign n20655_o = n20654_o[207];
  /* loadstore1.vhdl:708:59  */
  assign n20656_o = r2[299];
  /* loadstore1.vhdl:708:42  */
  assign n20657_o = ~n20656_o;
  /* loadstore1.vhdl:708:40  */
  assign n20659_o = {1'b1, n20657_o};
  /* loadstore1.vhdl:707:17  */
  assign n20661_o = n20655_o ? n20659_o : 2'b10;
  /* loadstore1.vhdl:706:13  */
  assign n20663_o = n20653_o ? n20661_o : 2'b00;
  /* loadstore1.vhdl:706:43  */
  assign n20664_o = r2[272:0];
  /* loadstore1.vhdl:706:47  */
  assign n20665_o = n20664_o[171:168];
  /* loadstore1.vhdl:706:20  */
  assign n20666_o = {27'b0, n20665_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20667_o = {1'b0, n20666_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20669_o = $signed(32'b00000000000000000000000000000011) < $signed(n20667_o);
  /* loadstore1.vhdl:707:23  */
  assign n20670_o = r2[272:0];
  /* loadstore1.vhdl:707:27  */
  assign n20671_o = n20670_o[207];
  /* loadstore1.vhdl:708:59  */
  assign n20672_o = r2[300];
  /* loadstore1.vhdl:708:42  */
  assign n20673_o = ~n20672_o;
  /* loadstore1.vhdl:708:40  */
  assign n20675_o = {1'b1, n20673_o};
  /* loadstore1.vhdl:707:17  */
  assign n20677_o = n20671_o ? n20675_o : 2'b10;
  /* loadstore1.vhdl:706:13  */
  assign n20679_o = n20669_o ? n20677_o : 2'b00;
  /* loadstore1.vhdl:706:43  */
  assign n20680_o = r2[272:0];
  /* loadstore1.vhdl:706:47  */
  assign n20681_o = n20680_o[171:168];
  /* loadstore1.vhdl:706:20  */
  assign n20682_o = {27'b0, n20681_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20683_o = {1'b0, n20682_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20685_o = $signed(32'b00000000000000000000000000000100) < $signed(n20683_o);
  /* loadstore1.vhdl:707:23  */
  assign n20686_o = r2[272:0];
  /* loadstore1.vhdl:707:27  */
  assign n20687_o = n20686_o[207];
  /* loadstore1.vhdl:708:59  */
  assign n20688_o = r2[301];
  /* loadstore1.vhdl:708:42  */
  assign n20689_o = ~n20688_o;
  /* loadstore1.vhdl:708:40  */
  assign n20691_o = {1'b1, n20689_o};
  /* loadstore1.vhdl:707:17  */
  assign n20693_o = n20687_o ? n20691_o : 2'b10;
  /* loadstore1.vhdl:706:13  */
  assign n20695_o = n20685_o ? n20693_o : 2'b00;
  /* loadstore1.vhdl:706:43  */
  assign n20696_o = r2[272:0];
  /* loadstore1.vhdl:706:47  */
  assign n20697_o = n20696_o[171:168];
  /* loadstore1.vhdl:706:20  */
  assign n20698_o = {27'b0, n20697_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20699_o = {1'b0, n20698_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20701_o = $signed(32'b00000000000000000000000000000101) < $signed(n20699_o);
  /* loadstore1.vhdl:707:23  */
  assign n20702_o = r2[272:0];
  /* loadstore1.vhdl:707:27  */
  assign n20703_o = n20702_o[207];
  /* loadstore1.vhdl:708:59  */
  assign n20704_o = r2[302];
  /* loadstore1.vhdl:708:42  */
  assign n20705_o = ~n20704_o;
  /* loadstore1.vhdl:708:40  */
  assign n20707_o = {1'b1, n20705_o};
  /* loadstore1.vhdl:707:17  */
  assign n20709_o = n20703_o ? n20707_o : 2'b10;
  /* loadstore1.vhdl:706:13  */
  assign n20711_o = n20701_o ? n20709_o : 2'b00;
  /* loadstore1.vhdl:706:43  */
  assign n20712_o = r2[272:0];
  /* loadstore1.vhdl:706:47  */
  assign n20713_o = n20712_o[171:168];
  /* loadstore1.vhdl:706:20  */
  assign n20714_o = {27'b0, n20713_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20715_o = {1'b0, n20714_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20717_o = $signed(32'b00000000000000000000000000000110) < $signed(n20715_o);
  /* loadstore1.vhdl:707:23  */
  assign n20718_o = r2[272:0];
  /* loadstore1.vhdl:707:27  */
  assign n20719_o = n20718_o[207];
  /* loadstore1.vhdl:708:59  */
  assign n20720_o = r2[303];
  /* loadstore1.vhdl:708:42  */
  assign n20721_o = ~n20720_o;
  /* loadstore1.vhdl:708:40  */
  assign n20723_o = {1'b1, n20721_o};
  /* loadstore1.vhdl:707:17  */
  assign n20725_o = n20719_o ? n20723_o : 2'b10;
  /* loadstore1.vhdl:706:13  */
  assign n20727_o = n20717_o ? n20725_o : 2'b00;
  /* loadstore1.vhdl:706:43  */
  assign n20728_o = r2[272:0];
  /* loadstore1.vhdl:706:47  */
  assign n20729_o = n20728_o[171:168];
  /* loadstore1.vhdl:706:20  */
  assign n20730_o = {27'b0, n20729_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20731_o = {1'b0, n20730_o};  //  uext
  /* loadstore1.vhdl:706:18  */
  assign n20733_o = $signed(32'b00000000000000000000000000000111) < $signed(n20731_o);
  /* loadstore1.vhdl:707:23  */
  assign n20734_o = r2[272:0];
  /* loadstore1.vhdl:707:27  */
  assign n20735_o = n20734_o[207];
  /* loadstore1.vhdl:708:59  */
  assign n20736_o = r2[304];
  /* loadstore1.vhdl:708:42  */
  assign n20737_o = ~n20736_o;
  /* loadstore1.vhdl:708:40  */
  assign n20739_o = {1'b1, n20737_o};
  /* loadstore1.vhdl:707:17  */
  assign n20741_o = n20735_o ? n20739_o : 2'b10;
  /* loadstore1.vhdl:706:13  */
  assign n20743_o = n20733_o ? n20741_o : 2'b00;
  assign n20744_o = {n20631_o, n20647_o, n20663_o, n20679_o, n20695_o, n20711_o, n20727_o, n20743_o};
  /* loadstore1.vhdl:718:26  */
  assign n20745_o = n20744_o[15:14];
  /* loadstore1.vhdl:720:73  */
  assign n20746_o = r3[92:85];
  /* loadstore1.vhdl:719:17  */
  assign n20748_o = n20745_o == 2'b11;
  assign n20749_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:722:74  */
  assign n20750_o = n20749_o[7:0];
  /* loadstore1.vhdl:721:17  */
  assign n20752_o = n20745_o == 2'b10;
  /* loadstore1.vhdl:724:88  */
  assign n20753_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20754_o = n20753_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20755_o = n20615_o & n20754_o;
  /* loadstore1.vhdl:724:88  */
  assign n20756_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20757_o = n20756_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20758_o = n20615_o & n20757_o;
  /* loadstore1.vhdl:724:88  */
  assign n20759_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20760_o = n20759_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20761_o = n20615_o & n20760_o;
  /* loadstore1.vhdl:724:88  */
  assign n20762_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20763_o = n20762_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20764_o = n20615_o & n20763_o;
  /* loadstore1.vhdl:724:88  */
  assign n20765_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20766_o = n20765_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20767_o = n20615_o & n20766_o;
  /* loadstore1.vhdl:724:88  */
  assign n20768_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20769_o = n20768_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20770_o = n20615_o & n20769_o;
  /* loadstore1.vhdl:724:88  */
  assign n20771_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20772_o = n20771_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20773_o = n20615_o & n20772_o;
  /* loadstore1.vhdl:724:88  */
  assign n20774_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20775_o = n20774_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20776_o = n20615_o & n20775_o;
  assign n20777_o = {n20755_o, n20758_o, n20761_o, n20764_o};
  assign n20778_o = {n20767_o, n20770_o, n20773_o, n20776_o};
  assign n20779_o = {n20777_o, n20778_o};
  assign n20780_o = {n20752_o, n20748_o};
  /* loadstore1.vhdl:718:13  */
  always @*
    case (n20780_o)
      2'b10: n20781_o = n20750_o;
      2'b01: n20781_o = n20746_o;
      default: n20781_o = n20779_o;
    endcase
  assign n20782_o = {n20631_o, n20647_o, n20663_o, n20679_o, n20695_o, n20711_o, n20727_o, n20743_o};
  /* loadstore1.vhdl:718:26  */
  assign n20783_o = n20782_o[13:12];
  /* loadstore1.vhdl:720:73  */
  assign n20784_o = r3[100:93];
  /* loadstore1.vhdl:719:17  */
  assign n20786_o = n20783_o == 2'b11;
  assign n20787_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:722:74  */
  assign n20788_o = n20787_o[15:8];
  /* loadstore1.vhdl:721:17  */
  assign n20790_o = n20783_o == 2'b10;
  /* loadstore1.vhdl:724:88  */
  assign n20791_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20792_o = n20791_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20793_o = n20615_o & n20792_o;
  /* loadstore1.vhdl:724:88  */
  assign n20794_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20795_o = n20794_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20796_o = n20615_o & n20795_o;
  /* loadstore1.vhdl:724:88  */
  assign n20797_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20798_o = n20797_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20799_o = n20615_o & n20798_o;
  /* loadstore1.vhdl:724:88  */
  assign n20800_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20801_o = n20800_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20802_o = n20615_o & n20801_o;
  /* loadstore1.vhdl:724:88  */
  assign n20803_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20804_o = n20803_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20805_o = n20615_o & n20804_o;
  /* loadstore1.vhdl:724:88  */
  assign n20806_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20807_o = n20806_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20808_o = n20615_o & n20807_o;
  /* loadstore1.vhdl:724:88  */
  assign n20809_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20810_o = n20809_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20811_o = n20615_o & n20810_o;
  /* loadstore1.vhdl:724:88  */
  assign n20812_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20813_o = n20812_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20814_o = n20615_o & n20813_o;
  assign n20815_o = {n20793_o, n20796_o, n20799_o, n20802_o};
  assign n20816_o = {n20805_o, n20808_o, n20811_o, n20814_o};
  assign n20817_o = {n20815_o, n20816_o};
  assign n20818_o = {n20790_o, n20786_o};
  /* loadstore1.vhdl:718:13  */
  always @*
    case (n20818_o)
      2'b10: n20819_o = n20788_o;
      2'b01: n20819_o = n20784_o;
      default: n20819_o = n20817_o;
    endcase
  assign n20820_o = {n20631_o, n20647_o, n20663_o, n20679_o, n20695_o, n20711_o, n20727_o, n20743_o};
  /* loadstore1.vhdl:718:26  */
  assign n20821_o = n20820_o[11:10];
  /* loadstore1.vhdl:720:73  */
  assign n20822_o = r3[108:101];
  /* loadstore1.vhdl:719:17  */
  assign n20824_o = n20821_o == 2'b11;
  assign n20825_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:722:74  */
  assign n20826_o = n20825_o[23:16];
  /* loadstore1.vhdl:721:17  */
  assign n20828_o = n20821_o == 2'b10;
  /* loadstore1.vhdl:724:88  */
  assign n20829_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20830_o = n20829_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20831_o = n20615_o & n20830_o;
  /* loadstore1.vhdl:724:88  */
  assign n20832_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20833_o = n20832_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20834_o = n20615_o & n20833_o;
  /* loadstore1.vhdl:724:88  */
  assign n20835_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20836_o = n20835_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20837_o = n20615_o & n20836_o;
  /* loadstore1.vhdl:724:88  */
  assign n20838_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20839_o = n20838_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20840_o = n20615_o & n20839_o;
  /* loadstore1.vhdl:724:88  */
  assign n20841_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20842_o = n20841_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20843_o = n20615_o & n20842_o;
  /* loadstore1.vhdl:724:88  */
  assign n20844_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20845_o = n20844_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20846_o = n20615_o & n20845_o;
  /* loadstore1.vhdl:724:88  */
  assign n20847_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20848_o = n20847_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20849_o = n20615_o & n20848_o;
  /* loadstore1.vhdl:724:88  */
  assign n20850_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20851_o = n20850_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20852_o = n20615_o & n20851_o;
  assign n20853_o = {n20831_o, n20834_o, n20837_o, n20840_o};
  assign n20854_o = {n20843_o, n20846_o, n20849_o, n20852_o};
  assign n20855_o = {n20853_o, n20854_o};
  assign n20856_o = {n20828_o, n20824_o};
  /* loadstore1.vhdl:718:13  */
  always @*
    case (n20856_o)
      2'b10: n20857_o = n20826_o;
      2'b01: n20857_o = n20822_o;
      default: n20857_o = n20855_o;
    endcase
  assign n20858_o = {n20631_o, n20647_o, n20663_o, n20679_o, n20695_o, n20711_o, n20727_o, n20743_o};
  /* loadstore1.vhdl:718:26  */
  assign n20859_o = n20858_o[9:8];
  /* loadstore1.vhdl:720:73  */
  assign n20860_o = r3[116:109];
  /* loadstore1.vhdl:719:17  */
  assign n20862_o = n20859_o == 2'b11;
  assign n20863_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:722:74  */
  assign n20864_o = n20863_o[31:24];
  /* loadstore1.vhdl:721:17  */
  assign n20866_o = n20859_o == 2'b10;
  /* loadstore1.vhdl:724:88  */
  assign n20867_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20868_o = n20867_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20869_o = n20615_o & n20868_o;
  /* loadstore1.vhdl:724:88  */
  assign n20870_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20871_o = n20870_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20872_o = n20615_o & n20871_o;
  /* loadstore1.vhdl:724:88  */
  assign n20873_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20874_o = n20873_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20875_o = n20615_o & n20874_o;
  /* loadstore1.vhdl:724:88  */
  assign n20876_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20877_o = n20876_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20878_o = n20615_o & n20877_o;
  /* loadstore1.vhdl:724:88  */
  assign n20879_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20880_o = n20879_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20881_o = n20615_o & n20880_o;
  /* loadstore1.vhdl:724:88  */
  assign n20882_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20883_o = n20882_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20884_o = n20615_o & n20883_o;
  /* loadstore1.vhdl:724:88  */
  assign n20885_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20886_o = n20885_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20887_o = n20615_o & n20886_o;
  /* loadstore1.vhdl:724:88  */
  assign n20888_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20889_o = n20888_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20890_o = n20615_o & n20889_o;
  assign n20891_o = {n20869_o, n20872_o, n20875_o, n20878_o};
  assign n20892_o = {n20881_o, n20884_o, n20887_o, n20890_o};
  assign n20893_o = {n20891_o, n20892_o};
  assign n20894_o = {n20866_o, n20862_o};
  /* loadstore1.vhdl:718:13  */
  always @*
    case (n20894_o)
      2'b10: n20895_o = n20864_o;
      2'b01: n20895_o = n20860_o;
      default: n20895_o = n20893_o;
    endcase
  assign n20896_o = {n20631_o, n20647_o, n20663_o, n20679_o, n20695_o, n20711_o, n20727_o, n20743_o};
  /* loadstore1.vhdl:718:26  */
  assign n20897_o = n20896_o[7:6];
  /* loadstore1.vhdl:720:73  */
  assign n20898_o = r3[124:117];
  /* loadstore1.vhdl:719:17  */
  assign n20900_o = n20897_o == 2'b11;
  assign n20901_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:722:74  */
  assign n20902_o = n20901_o[39:32];
  /* loadstore1.vhdl:721:17  */
  assign n20904_o = n20897_o == 2'b10;
  /* loadstore1.vhdl:724:88  */
  assign n20905_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20906_o = n20905_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20907_o = n20615_o & n20906_o;
  /* loadstore1.vhdl:724:88  */
  assign n20908_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20909_o = n20908_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20910_o = n20615_o & n20909_o;
  /* loadstore1.vhdl:724:88  */
  assign n20911_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20912_o = n20911_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20913_o = n20615_o & n20912_o;
  /* loadstore1.vhdl:724:88  */
  assign n20914_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20915_o = n20914_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20916_o = n20615_o & n20915_o;
  /* loadstore1.vhdl:724:88  */
  assign n20917_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20918_o = n20917_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20919_o = n20615_o & n20918_o;
  /* loadstore1.vhdl:724:88  */
  assign n20920_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20921_o = n20920_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20922_o = n20615_o & n20921_o;
  /* loadstore1.vhdl:724:88  */
  assign n20923_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20924_o = n20923_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20925_o = n20615_o & n20924_o;
  /* loadstore1.vhdl:724:88  */
  assign n20926_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20927_o = n20926_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20928_o = n20615_o & n20927_o;
  assign n20929_o = {n20907_o, n20910_o, n20913_o, n20916_o};
  assign n20930_o = {n20919_o, n20922_o, n20925_o, n20928_o};
  assign n20931_o = {n20929_o, n20930_o};
  assign n20932_o = {n20904_o, n20900_o};
  /* loadstore1.vhdl:718:13  */
  always @*
    case (n20932_o)
      2'b10: n20933_o = n20902_o;
      2'b01: n20933_o = n20898_o;
      default: n20933_o = n20931_o;
    endcase
  assign n20934_o = {n20631_o, n20647_o, n20663_o, n20679_o, n20695_o, n20711_o, n20727_o, n20743_o};
  /* loadstore1.vhdl:718:26  */
  assign n20935_o = n20934_o[5:4];
  /* loadstore1.vhdl:720:73  */
  assign n20936_o = r3[132:125];
  /* loadstore1.vhdl:719:17  */
  assign n20938_o = n20935_o == 2'b11;
  assign n20939_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:722:74  */
  assign n20940_o = n20939_o[47:40];
  /* loadstore1.vhdl:721:17  */
  assign n20942_o = n20935_o == 2'b10;
  /* loadstore1.vhdl:724:88  */
  assign n20943_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20944_o = n20943_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20945_o = n20615_o & n20944_o;
  /* loadstore1.vhdl:724:88  */
  assign n20946_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20947_o = n20946_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20948_o = n20615_o & n20947_o;
  /* loadstore1.vhdl:724:88  */
  assign n20949_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20950_o = n20949_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20951_o = n20615_o & n20950_o;
  /* loadstore1.vhdl:724:88  */
  assign n20952_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20953_o = n20952_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20954_o = n20615_o & n20953_o;
  /* loadstore1.vhdl:724:88  */
  assign n20955_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20956_o = n20955_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20957_o = n20615_o & n20956_o;
  /* loadstore1.vhdl:724:88  */
  assign n20958_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20959_o = n20958_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20960_o = n20615_o & n20959_o;
  /* loadstore1.vhdl:724:88  */
  assign n20961_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20962_o = n20961_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20963_o = n20615_o & n20962_o;
  /* loadstore1.vhdl:724:88  */
  assign n20964_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20965_o = n20964_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20966_o = n20615_o & n20965_o;
  assign n20967_o = {n20945_o, n20948_o, n20951_o, n20954_o};
  assign n20968_o = {n20957_o, n20960_o, n20963_o, n20966_o};
  assign n20969_o = {n20967_o, n20968_o};
  assign n20970_o = {n20942_o, n20938_o};
  /* loadstore1.vhdl:718:13  */
  always @*
    case (n20970_o)
      2'b10: n20971_o = n20940_o;
      2'b01: n20971_o = n20936_o;
      default: n20971_o = n20969_o;
    endcase
  assign n20972_o = {n20631_o, n20647_o, n20663_o, n20679_o, n20695_o, n20711_o, n20727_o, n20743_o};
  /* loadstore1.vhdl:718:26  */
  assign n20973_o = n20972_o[3:2];
  /* loadstore1.vhdl:720:73  */
  assign n20974_o = r3[140:133];
  /* loadstore1.vhdl:719:17  */
  assign n20976_o = n20973_o == 2'b11;
  assign n20977_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:722:74  */
  assign n20978_o = n20977_o[55:48];
  /* loadstore1.vhdl:721:17  */
  assign n20980_o = n20973_o == 2'b10;
  /* loadstore1.vhdl:724:88  */
  assign n20981_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20982_o = n20981_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20983_o = n20615_o & n20982_o;
  /* loadstore1.vhdl:724:88  */
  assign n20984_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20985_o = n20984_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20986_o = n20615_o & n20985_o;
  /* loadstore1.vhdl:724:88  */
  assign n20987_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20988_o = n20987_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20989_o = n20615_o & n20988_o;
  /* loadstore1.vhdl:724:88  */
  assign n20990_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20991_o = n20990_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20992_o = n20615_o & n20991_o;
  /* loadstore1.vhdl:724:88  */
  assign n20993_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20994_o = n20993_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20995_o = n20615_o & n20994_o;
  /* loadstore1.vhdl:724:88  */
  assign n20996_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n20997_o = n20996_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n20998_o = n20615_o & n20997_o;
  /* loadstore1.vhdl:724:88  */
  assign n20999_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n21000_o = n20999_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n21001_o = n20615_o & n21000_o;
  /* loadstore1.vhdl:724:88  */
  assign n21002_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n21003_o = n21002_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n21004_o = n20615_o & n21003_o;
  assign n21005_o = {n20983_o, n20986_o, n20989_o, n20992_o};
  assign n21006_o = {n20995_o, n20998_o, n21001_o, n21004_o};
  assign n21007_o = {n21005_o, n21006_o};
  assign n21008_o = {n20980_o, n20976_o};
  /* loadstore1.vhdl:718:13  */
  always @*
    case (n21008_o)
      2'b10: n21009_o = n20978_o;
      2'b01: n21009_o = n20974_o;
      default: n21009_o = n21007_o;
    endcase
  assign n21010_o = {n20631_o, n20647_o, n20663_o, n20679_o, n20695_o, n20711_o, n20727_o, n20743_o};
  /* loadstore1.vhdl:718:26  */
  assign n21011_o = n21010_o[1:0];
  /* loadstore1.vhdl:720:73  */
  assign n21012_o = r3[148:141];
  /* loadstore1.vhdl:719:17  */
  assign n21014_o = n21011_o == 2'b11;
  assign n21015_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  /* loadstore1.vhdl:722:74  */
  assign n21016_o = n21015_o[63:56];
  /* loadstore1.vhdl:721:17  */
  assign n21018_o = n21011_o == 2'b10;
  /* loadstore1.vhdl:724:88  */
  assign n21019_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n21020_o = n21019_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n21021_o = n20615_o & n21020_o;
  /* loadstore1.vhdl:724:88  */
  assign n21022_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n21023_o = n21022_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n21024_o = n20615_o & n21023_o;
  /* loadstore1.vhdl:724:88  */
  assign n21025_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n21026_o = n21025_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n21027_o = n20615_o & n21026_o;
  /* loadstore1.vhdl:724:88  */
  assign n21028_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n21029_o = n21028_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n21030_o = n20615_o & n21029_o;
  /* loadstore1.vhdl:724:88  */
  assign n21031_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n21032_o = n21031_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n21033_o = n20615_o & n21032_o;
  /* loadstore1.vhdl:724:88  */
  assign n21034_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n21035_o = n21034_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n21036_o = n20615_o & n21035_o;
  /* loadstore1.vhdl:724:88  */
  assign n21037_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n21038_o = n21037_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n21039_o = n20615_o & n21038_o;
  /* loadstore1.vhdl:724:88  */
  assign n21040_o = r2[272:0];
  /* loadstore1.vhdl:724:92  */
  assign n21041_o = n21040_o[180];
  /* loadstore1.vhdl:724:81  */
  assign n21042_o = n20615_o & n21041_o;
  assign n21043_o = {n21021_o, n21024_o, n21027_o, n21030_o};
  assign n21044_o = {n21033_o, n21036_o, n21039_o, n21042_o};
  assign n21045_o = {n21043_o, n21044_o};
  assign n21046_o = {n21018_o, n21014_o};
  /* loadstore1.vhdl:718:13  */
  always @*
    case (n21046_o)
      2'b10: n21047_o = n21016_o;
      2'b01: n21047_o = n21012_o;
      default: n21047_o = n21045_o;
    endcase
  assign n21048_o = {n21047_o, n21009_o, n20971_o, n20933_o, n20895_o, n20857_o, n20819_o, n20781_o};
  /* loadstore1.vhdl:730:41  */
  assign n21049_o = n21048_o[31:0];
  assign n21052_o = {n21047_o, n21009_o, n20971_o, n20933_o, n20895_o, n20857_o, n20819_o, n20781_o};
  /* loadstore1.vhdl:731:43  */
  assign n21053_o = n21052_o[22:0];
  /* loadstore1.vhdl:731:27  */
  assign n21054_o = |(n21053_o);
  assign n21057_o = {n21047_o, n21009_o, n20971_o, n20933_o, n20895_o, n20857_o, n20819_o, n20781_o};
  /* loadstore1.vhdl:732:57  */
  assign n21058_o = n21057_o[22:0];
  /* helpers.vhdl:221:43  */
  assign n21070_o = n21058_o[0];
  /* helpers.vhdl:221:43  */
  assign n21073_o = n21058_o[1];
  /* helpers.vhdl:221:43  */
  assign n21075_o = n21058_o[2];
  /* helpers.vhdl:221:43  */
  assign n21077_o = n21058_o[3];
  /* helpers.vhdl:221:43  */
  assign n21079_o = n21058_o[4];
  /* helpers.vhdl:221:43  */
  assign n21081_o = n21058_o[5];
  /* helpers.vhdl:221:43  */
  assign n21083_o = n21058_o[6];
  /* helpers.vhdl:221:43  */
  assign n21085_o = n21058_o[7];
  /* helpers.vhdl:221:43  */
  assign n21087_o = n21058_o[8];
  /* helpers.vhdl:221:43  */
  assign n21089_o = n21058_o[9];
  /* helpers.vhdl:221:43  */
  assign n21091_o = n21058_o[10];
  /* helpers.vhdl:221:43  */
  assign n21093_o = n21058_o[11];
  /* helpers.vhdl:221:43  */
  assign n21095_o = n21058_o[12];
  /* helpers.vhdl:221:43  */
  assign n21097_o = n21058_o[13];
  /* helpers.vhdl:221:43  */
  assign n21099_o = n21058_o[14];
  /* helpers.vhdl:221:43  */
  assign n21101_o = n21058_o[15];
  /* helpers.vhdl:221:43  */
  assign n21103_o = n21058_o[16];
  /* helpers.vhdl:221:43  */
  assign n21105_o = n21058_o[17];
  /* helpers.vhdl:221:43  */
  assign n21107_o = n21058_o[18];
  /* helpers.vhdl:221:43  */
  assign n21109_o = n21058_o[19];
  /* helpers.vhdl:221:43  */
  assign n21111_o = n21058_o[20];
  /* helpers.vhdl:221:43  */
  assign n21113_o = n21058_o[21];
  /* helpers.vhdl:221:43  */
  assign n21115_o = n21058_o[22];
  assign n21116_o = {n21070_o, n21073_o, n21075_o, n21077_o, n21079_o, n21081_o, n21083_o, n21085_o, n21087_o, n21089_o, n21091_o, n21093_o, n21095_o, n21097_o, n21099_o, n21101_o, n21103_o, n21105_o, n21107_o, n21109_o, n21111_o, n21113_o, n21115_o};
  /* helpers.vhdl:282:34  */
  assign n21129_o = -n21116_o;
  /* helpers.vhdl:283:23  */
  assign n21131_o = n21129_o & n21116_o;
  /* helpers.vhdl:284:21  */
  assign n21133_o = n21129_o | n21116_o;
  /* helpers.vhdl:285:48  */
  assign n21136_o = {{41{n21133_o[22]}}, n21133_o}; // sext
  /* helpers.vhdl:266:29  */
  assign n21145_o = n21136_o[1];
  /* helpers.vhdl:266:55  */
  assign n21146_o = n21136_o[0];
  /* helpers.vhdl:266:50  */
  assign n21147_o = ~n21146_o;
  /* helpers.vhdl:266:46  */
  assign n21148_o = n21145_o & n21147_o;
  /* helpers.vhdl:266:24  */
  assign n21150_o = 1'b0 | n21148_o;
  /* helpers.vhdl:266:29  */
  assign n21152_o = n21136_o[3];
  /* helpers.vhdl:266:55  */
  assign n21153_o = n21136_o[2];
  /* helpers.vhdl:266:50  */
  assign n21154_o = ~n21153_o;
  /* helpers.vhdl:266:46  */
  assign n21155_o = n21152_o & n21154_o;
  /* helpers.vhdl:266:24  */
  assign n21156_o = n21150_o | n21155_o;
  /* helpers.vhdl:266:29  */
  assign n21157_o = n21136_o[5];
  /* helpers.vhdl:266:55  */
  assign n21158_o = n21136_o[4];
  /* helpers.vhdl:266:50  */
  assign n21159_o = ~n21158_o;
  /* helpers.vhdl:266:46  */
  assign n21160_o = n21157_o & n21159_o;
  /* helpers.vhdl:266:24  */
  assign n21161_o = n21156_o | n21160_o;
  /* helpers.vhdl:266:29  */
  assign n21162_o = n21136_o[7];
  /* helpers.vhdl:266:55  */
  assign n21163_o = n21136_o[6];
  /* helpers.vhdl:266:50  */
  assign n21164_o = ~n21163_o;
  /* helpers.vhdl:266:46  */
  assign n21165_o = n21162_o & n21164_o;
  /* helpers.vhdl:266:24  */
  assign n21166_o = n21161_o | n21165_o;
  /* helpers.vhdl:266:29  */
  assign n21167_o = n21136_o[9];
  /* helpers.vhdl:266:55  */
  assign n21168_o = n21136_o[8];
  /* helpers.vhdl:266:50  */
  assign n21169_o = ~n21168_o;
  /* helpers.vhdl:266:46  */
  assign n21170_o = n21167_o & n21169_o;
  /* helpers.vhdl:266:24  */
  assign n21171_o = n21166_o | n21170_o;
  /* helpers.vhdl:266:29  */
  assign n21172_o = n21136_o[11];
  /* helpers.vhdl:266:55  */
  assign n21173_o = n21136_o[10];
  /* helpers.vhdl:266:50  */
  assign n21174_o = ~n21173_o;
  /* helpers.vhdl:266:46  */
  assign n21175_o = n21172_o & n21174_o;
  /* helpers.vhdl:266:24  */
  assign n21176_o = n21171_o | n21175_o;
  /* helpers.vhdl:266:29  */
  assign n21177_o = n21136_o[13];
  /* helpers.vhdl:266:55  */
  assign n21178_o = n21136_o[12];
  /* helpers.vhdl:266:50  */
  assign n21179_o = ~n21178_o;
  /* helpers.vhdl:266:46  */
  assign n21180_o = n21177_o & n21179_o;
  /* helpers.vhdl:266:24  */
  assign n21181_o = n21176_o | n21180_o;
  /* helpers.vhdl:266:29  */
  assign n21182_o = n21136_o[15];
  /* helpers.vhdl:266:55  */
  assign n21183_o = n21136_o[14];
  /* helpers.vhdl:266:50  */
  assign n21184_o = ~n21183_o;
  /* helpers.vhdl:266:46  */
  assign n21185_o = n21182_o & n21184_o;
  /* helpers.vhdl:266:24  */
  assign n21186_o = n21181_o | n21185_o;
  /* helpers.vhdl:266:29  */
  assign n21187_o = n21136_o[17];
  /* helpers.vhdl:266:55  */
  assign n21188_o = n21136_o[16];
  /* helpers.vhdl:266:50  */
  assign n21189_o = ~n21188_o;
  /* helpers.vhdl:266:46  */
  assign n21190_o = n21187_o & n21189_o;
  /* helpers.vhdl:266:24  */
  assign n21191_o = n21186_o | n21190_o;
  /* helpers.vhdl:266:29  */
  assign n21192_o = n21136_o[19];
  /* helpers.vhdl:266:55  */
  assign n21193_o = n21136_o[18];
  /* helpers.vhdl:266:50  */
  assign n21194_o = ~n21193_o;
  /* helpers.vhdl:266:46  */
  assign n21195_o = n21192_o & n21194_o;
  /* helpers.vhdl:266:24  */
  assign n21196_o = n21191_o | n21195_o;
  /* helpers.vhdl:266:29  */
  assign n21197_o = n21136_o[21];
  /* helpers.vhdl:266:55  */
  assign n21198_o = n21136_o[20];
  /* helpers.vhdl:266:50  */
  assign n21199_o = ~n21198_o;
  /* helpers.vhdl:266:46  */
  assign n21200_o = n21197_o & n21199_o;
  /* helpers.vhdl:266:24  */
  assign n21201_o = n21196_o | n21200_o;
  /* helpers.vhdl:266:29  */
  assign n21202_o = n21136_o[23];
  /* helpers.vhdl:266:55  */
  assign n21203_o = n21136_o[22];
  /* helpers.vhdl:266:50  */
  assign n21204_o = ~n21203_o;
  /* helpers.vhdl:266:46  */
  assign n21205_o = n21202_o & n21204_o;
  /* helpers.vhdl:266:24  */
  assign n21206_o = n21201_o | n21205_o;
  /* helpers.vhdl:266:29  */
  assign n21207_o = n21136_o[25];
  /* helpers.vhdl:266:55  */
  assign n21208_o = n21136_o[24];
  /* helpers.vhdl:266:50  */
  assign n21209_o = ~n21208_o;
  /* helpers.vhdl:266:46  */
  assign n21210_o = n21207_o & n21209_o;
  /* helpers.vhdl:266:24  */
  assign n21211_o = n21206_o | n21210_o;
  /* helpers.vhdl:266:29  */
  assign n21212_o = n21136_o[27];
  /* helpers.vhdl:266:55  */
  assign n21213_o = n21136_o[26];
  /* helpers.vhdl:266:50  */
  assign n21214_o = ~n21213_o;
  /* helpers.vhdl:266:46  */
  assign n21215_o = n21212_o & n21214_o;
  /* helpers.vhdl:266:24  */
  assign n21216_o = n21211_o | n21215_o;
  /* helpers.vhdl:266:29  */
  assign n21217_o = n21136_o[29];
  /* helpers.vhdl:266:55  */
  assign n21218_o = n21136_o[28];
  /* helpers.vhdl:266:50  */
  assign n21219_o = ~n21218_o;
  /* helpers.vhdl:266:46  */
  assign n21220_o = n21217_o & n21219_o;
  /* helpers.vhdl:266:24  */
  assign n21221_o = n21216_o | n21220_o;
  /* helpers.vhdl:266:29  */
  assign n21222_o = n21136_o[31];
  /* helpers.vhdl:266:55  */
  assign n21223_o = n21136_o[30];
  /* helpers.vhdl:266:50  */
  assign n21224_o = ~n21223_o;
  /* helpers.vhdl:266:46  */
  assign n21225_o = n21222_o & n21224_o;
  /* helpers.vhdl:266:24  */
  assign n21226_o = n21221_o | n21225_o;
  /* helpers.vhdl:266:29  */
  assign n21227_o = n21136_o[33];
  /* helpers.vhdl:266:55  */
  assign n21228_o = n21136_o[32];
  /* helpers.vhdl:266:50  */
  assign n21229_o = ~n21228_o;
  /* helpers.vhdl:266:46  */
  assign n21230_o = n21227_o & n21229_o;
  /* helpers.vhdl:266:24  */
  assign n21231_o = n21226_o | n21230_o;
  /* helpers.vhdl:266:29  */
  assign n21232_o = n21136_o[35];
  /* helpers.vhdl:266:55  */
  assign n21233_o = n21136_o[34];
  /* helpers.vhdl:266:50  */
  assign n21234_o = ~n21233_o;
  /* helpers.vhdl:266:46  */
  assign n21235_o = n21232_o & n21234_o;
  /* helpers.vhdl:266:24  */
  assign n21236_o = n21231_o | n21235_o;
  /* helpers.vhdl:266:29  */
  assign n21237_o = n21136_o[37];
  /* helpers.vhdl:266:55  */
  assign n21238_o = n21136_o[36];
  /* helpers.vhdl:266:50  */
  assign n21239_o = ~n21238_o;
  /* helpers.vhdl:266:46  */
  assign n21240_o = n21237_o & n21239_o;
  /* helpers.vhdl:266:24  */
  assign n21241_o = n21236_o | n21240_o;
  /* helpers.vhdl:266:29  */
  assign n21242_o = n21136_o[39];
  /* helpers.vhdl:266:55  */
  assign n21243_o = n21136_o[38];
  /* helpers.vhdl:266:50  */
  assign n21244_o = ~n21243_o;
  /* helpers.vhdl:266:46  */
  assign n21245_o = n21242_o & n21244_o;
  /* helpers.vhdl:266:24  */
  assign n21246_o = n21241_o | n21245_o;
  /* helpers.vhdl:266:29  */
  assign n21247_o = n21136_o[41];
  /* helpers.vhdl:266:55  */
  assign n21248_o = n21136_o[40];
  /* helpers.vhdl:266:50  */
  assign n21249_o = ~n21248_o;
  /* helpers.vhdl:266:46  */
  assign n21250_o = n21247_o & n21249_o;
  /* helpers.vhdl:266:24  */
  assign n21251_o = n21246_o | n21250_o;
  /* helpers.vhdl:266:29  */
  assign n21252_o = n21136_o[43];
  /* helpers.vhdl:266:55  */
  assign n21253_o = n21136_o[42];
  /* helpers.vhdl:266:50  */
  assign n21254_o = ~n21253_o;
  /* helpers.vhdl:266:46  */
  assign n21255_o = n21252_o & n21254_o;
  /* helpers.vhdl:266:24  */
  assign n21256_o = n21251_o | n21255_o;
  /* helpers.vhdl:266:29  */
  assign n21257_o = n21136_o[45];
  /* helpers.vhdl:266:55  */
  assign n21258_o = n21136_o[44];
  /* helpers.vhdl:266:50  */
  assign n21259_o = ~n21258_o;
  /* helpers.vhdl:266:46  */
  assign n21260_o = n21257_o & n21259_o;
  /* helpers.vhdl:266:24  */
  assign n21261_o = n21256_o | n21260_o;
  /* helpers.vhdl:266:29  */
  assign n21262_o = n21136_o[47];
  /* helpers.vhdl:266:55  */
  assign n21263_o = n21136_o[46];
  /* helpers.vhdl:266:50  */
  assign n21264_o = ~n21263_o;
  /* helpers.vhdl:266:46  */
  assign n21265_o = n21262_o & n21264_o;
  /* helpers.vhdl:266:24  */
  assign n21266_o = n21261_o | n21265_o;
  /* helpers.vhdl:266:29  */
  assign n21267_o = n21136_o[49];
  /* helpers.vhdl:266:55  */
  assign n21268_o = n21136_o[48];
  /* helpers.vhdl:266:50  */
  assign n21269_o = ~n21268_o;
  /* helpers.vhdl:266:46  */
  assign n21270_o = n21267_o & n21269_o;
  /* helpers.vhdl:266:24  */
  assign n21271_o = n21266_o | n21270_o;
  /* helpers.vhdl:266:29  */
  assign n21272_o = n21136_o[51];
  /* helpers.vhdl:266:55  */
  assign n21273_o = n21136_o[50];
  /* helpers.vhdl:266:50  */
  assign n21274_o = ~n21273_o;
  /* helpers.vhdl:266:46  */
  assign n21275_o = n21272_o & n21274_o;
  /* helpers.vhdl:266:24  */
  assign n21276_o = n21271_o | n21275_o;
  /* helpers.vhdl:266:29  */
  assign n21277_o = n21136_o[53];
  /* helpers.vhdl:266:55  */
  assign n21278_o = n21136_o[52];
  /* helpers.vhdl:266:50  */
  assign n21279_o = ~n21278_o;
  /* helpers.vhdl:266:46  */
  assign n21280_o = n21277_o & n21279_o;
  /* helpers.vhdl:266:24  */
  assign n21281_o = n21276_o | n21280_o;
  /* helpers.vhdl:266:29  */
  assign n21282_o = n21136_o[55];
  /* helpers.vhdl:266:55  */
  assign n21283_o = n21136_o[54];
  /* helpers.vhdl:266:50  */
  assign n21284_o = ~n21283_o;
  /* helpers.vhdl:266:46  */
  assign n21285_o = n21282_o & n21284_o;
  /* helpers.vhdl:266:24  */
  assign n21286_o = n21281_o | n21285_o;
  /* helpers.vhdl:266:29  */
  assign n21287_o = n21136_o[57];
  /* helpers.vhdl:266:55  */
  assign n21288_o = n21136_o[56];
  /* helpers.vhdl:266:50  */
  assign n21289_o = ~n21288_o;
  /* helpers.vhdl:266:46  */
  assign n21290_o = n21287_o & n21289_o;
  /* helpers.vhdl:266:24  */
  assign n21291_o = n21286_o | n21290_o;
  /* helpers.vhdl:266:29  */
  assign n21292_o = n21136_o[59];
  /* helpers.vhdl:266:55  */
  assign n21293_o = n21136_o[58];
  /* helpers.vhdl:266:50  */
  assign n21294_o = ~n21293_o;
  /* helpers.vhdl:266:46  */
  assign n21295_o = n21292_o & n21294_o;
  /* helpers.vhdl:266:24  */
  assign n21296_o = n21291_o | n21295_o;
  /* helpers.vhdl:266:29  */
  assign n21297_o = n21136_o[61];
  /* helpers.vhdl:266:55  */
  assign n21298_o = n21136_o[60];
  /* helpers.vhdl:266:50  */
  assign n21299_o = ~n21298_o;
  /* helpers.vhdl:266:46  */
  assign n21300_o = n21297_o & n21299_o;
  /* helpers.vhdl:266:24  */
  assign n21301_o = n21296_o | n21300_o;
  /* helpers.vhdl:266:29  */
  assign n21302_o = n21136_o[63];
  /* helpers.vhdl:266:55  */
  assign n21303_o = n21136_o[62];
  /* helpers.vhdl:266:50  */
  assign n21304_o = ~n21303_o;
  /* helpers.vhdl:266:46  */
  assign n21305_o = n21302_o & n21304_o;
  /* helpers.vhdl:266:24  */
  assign n21306_o = n21301_o | n21305_o;
  /* helpers.vhdl:266:29  */
  assign n21309_o = n21136_o[3];
  /* helpers.vhdl:266:55  */
  assign n21310_o = n21136_o[1];
  /* helpers.vhdl:266:50  */
  assign n21311_o = ~n21310_o;
  /* helpers.vhdl:266:46  */
  assign n21312_o = n21309_o & n21311_o;
  /* helpers.vhdl:266:24  */
  assign n21314_o = 1'b0 | n21312_o;
  /* helpers.vhdl:266:29  */
  assign n21316_o = n21136_o[7];
  /* helpers.vhdl:266:55  */
  assign n21317_o = n21136_o[5];
  /* helpers.vhdl:266:50  */
  assign n21318_o = ~n21317_o;
  /* helpers.vhdl:266:46  */
  assign n21319_o = n21316_o & n21318_o;
  /* helpers.vhdl:266:24  */
  assign n21320_o = n21314_o | n21319_o;
  /* helpers.vhdl:266:29  */
  assign n21321_o = n21136_o[11];
  /* helpers.vhdl:266:55  */
  assign n21322_o = n21136_o[9];
  /* helpers.vhdl:266:50  */
  assign n21323_o = ~n21322_o;
  /* helpers.vhdl:266:46  */
  assign n21324_o = n21321_o & n21323_o;
  /* helpers.vhdl:266:24  */
  assign n21325_o = n21320_o | n21324_o;
  /* helpers.vhdl:266:29  */
  assign n21326_o = n21136_o[15];
  /* helpers.vhdl:266:55  */
  assign n21327_o = n21136_o[13];
  /* helpers.vhdl:266:50  */
  assign n21328_o = ~n21327_o;
  /* helpers.vhdl:266:46  */
  assign n21329_o = n21326_o & n21328_o;
  /* helpers.vhdl:266:24  */
  assign n21330_o = n21325_o | n21329_o;
  /* helpers.vhdl:266:29  */
  assign n21331_o = n21136_o[19];
  /* helpers.vhdl:266:55  */
  assign n21332_o = n21136_o[17];
  /* helpers.vhdl:266:50  */
  assign n21333_o = ~n21332_o;
  /* helpers.vhdl:266:46  */
  assign n21334_o = n21331_o & n21333_o;
  /* helpers.vhdl:266:24  */
  assign n21335_o = n21330_o | n21334_o;
  /* helpers.vhdl:266:29  */
  assign n21336_o = n21136_o[23];
  /* helpers.vhdl:266:55  */
  assign n21337_o = n21136_o[21];
  /* helpers.vhdl:266:50  */
  assign n21338_o = ~n21337_o;
  /* helpers.vhdl:266:46  */
  assign n21339_o = n21336_o & n21338_o;
  /* helpers.vhdl:266:24  */
  assign n21340_o = n21335_o | n21339_o;
  /* helpers.vhdl:266:29  */
  assign n21341_o = n21136_o[27];
  /* helpers.vhdl:266:55  */
  assign n21342_o = n21136_o[25];
  /* helpers.vhdl:266:50  */
  assign n21343_o = ~n21342_o;
  /* helpers.vhdl:266:46  */
  assign n21344_o = n21341_o & n21343_o;
  /* helpers.vhdl:266:24  */
  assign n21345_o = n21340_o | n21344_o;
  /* helpers.vhdl:266:29  */
  assign n21346_o = n21136_o[31];
  /* helpers.vhdl:266:55  */
  assign n21347_o = n21136_o[29];
  /* helpers.vhdl:266:50  */
  assign n21348_o = ~n21347_o;
  /* helpers.vhdl:266:46  */
  assign n21349_o = n21346_o & n21348_o;
  /* helpers.vhdl:266:24  */
  assign n21350_o = n21345_o | n21349_o;
  /* helpers.vhdl:266:29  */
  assign n21351_o = n21136_o[35];
  /* helpers.vhdl:266:55  */
  assign n21352_o = n21136_o[33];
  /* helpers.vhdl:266:50  */
  assign n21353_o = ~n21352_o;
  /* helpers.vhdl:266:46  */
  assign n21354_o = n21351_o & n21353_o;
  /* helpers.vhdl:266:24  */
  assign n21355_o = n21350_o | n21354_o;
  /* helpers.vhdl:266:29  */
  assign n21356_o = n21136_o[39];
  /* helpers.vhdl:266:55  */
  assign n21357_o = n21136_o[37];
  /* helpers.vhdl:266:50  */
  assign n21358_o = ~n21357_o;
  /* helpers.vhdl:266:46  */
  assign n21359_o = n21356_o & n21358_o;
  /* helpers.vhdl:266:24  */
  assign n21360_o = n21355_o | n21359_o;
  /* helpers.vhdl:266:29  */
  assign n21361_o = n21136_o[43];
  /* helpers.vhdl:266:55  */
  assign n21362_o = n21136_o[41];
  /* helpers.vhdl:266:50  */
  assign n21363_o = ~n21362_o;
  /* helpers.vhdl:266:46  */
  assign n21364_o = n21361_o & n21363_o;
  /* helpers.vhdl:266:24  */
  assign n21365_o = n21360_o | n21364_o;
  /* helpers.vhdl:266:29  */
  assign n21366_o = n21136_o[47];
  /* helpers.vhdl:266:55  */
  assign n21367_o = n21136_o[45];
  /* helpers.vhdl:266:50  */
  assign n21368_o = ~n21367_o;
  /* helpers.vhdl:266:46  */
  assign n21369_o = n21366_o & n21368_o;
  /* helpers.vhdl:266:24  */
  assign n21370_o = n21365_o | n21369_o;
  /* helpers.vhdl:266:29  */
  assign n21371_o = n21136_o[51];
  /* helpers.vhdl:266:55  */
  assign n21372_o = n21136_o[49];
  /* helpers.vhdl:266:50  */
  assign n21373_o = ~n21372_o;
  /* helpers.vhdl:266:46  */
  assign n21374_o = n21371_o & n21373_o;
  /* helpers.vhdl:266:24  */
  assign n21375_o = n21370_o | n21374_o;
  /* helpers.vhdl:266:29  */
  assign n21376_o = n21136_o[55];
  /* helpers.vhdl:266:55  */
  assign n21377_o = n21136_o[53];
  /* helpers.vhdl:266:50  */
  assign n21378_o = ~n21377_o;
  /* helpers.vhdl:266:46  */
  assign n21379_o = n21376_o & n21378_o;
  /* helpers.vhdl:266:24  */
  assign n21380_o = n21375_o | n21379_o;
  /* helpers.vhdl:266:29  */
  assign n21381_o = n21136_o[59];
  /* helpers.vhdl:266:55  */
  assign n21382_o = n21136_o[57];
  /* helpers.vhdl:266:50  */
  assign n21383_o = ~n21382_o;
  /* helpers.vhdl:266:46  */
  assign n21384_o = n21381_o & n21383_o;
  /* helpers.vhdl:266:24  */
  assign n21385_o = n21380_o | n21384_o;
  /* helpers.vhdl:266:29  */
  assign n21386_o = n21136_o[63];
  /* helpers.vhdl:266:55  */
  assign n21387_o = n21136_o[61];
  /* helpers.vhdl:266:50  */
  assign n21388_o = ~n21387_o;
  /* helpers.vhdl:266:46  */
  assign n21389_o = n21386_o & n21388_o;
  /* helpers.vhdl:266:24  */
  assign n21390_o = n21385_o | n21389_o;
  /* helpers.vhdl:266:29  */
  assign n21392_o = n21136_o[7];
  /* helpers.vhdl:266:55  */
  assign n21393_o = n21136_o[3];
  /* helpers.vhdl:266:50  */
  assign n21394_o = ~n21393_o;
  /* helpers.vhdl:266:46  */
  assign n21395_o = n21392_o & n21394_o;
  /* helpers.vhdl:266:24  */
  assign n21397_o = 1'b0 | n21395_o;
  /* helpers.vhdl:266:29  */
  assign n21399_o = n21136_o[15];
  /* helpers.vhdl:266:55  */
  assign n21400_o = n21136_o[11];
  /* helpers.vhdl:266:50  */
  assign n21401_o = ~n21400_o;
  /* helpers.vhdl:266:46  */
  assign n21402_o = n21399_o & n21401_o;
  /* helpers.vhdl:266:24  */
  assign n21403_o = n21397_o | n21402_o;
  /* helpers.vhdl:266:29  */
  assign n21404_o = n21136_o[23];
  /* helpers.vhdl:266:55  */
  assign n21405_o = n21136_o[19];
  /* helpers.vhdl:266:50  */
  assign n21406_o = ~n21405_o;
  /* helpers.vhdl:266:46  */
  assign n21407_o = n21404_o & n21406_o;
  /* helpers.vhdl:266:24  */
  assign n21408_o = n21403_o | n21407_o;
  /* helpers.vhdl:266:29  */
  assign n21409_o = n21136_o[31];
  /* helpers.vhdl:266:55  */
  assign n21410_o = n21136_o[27];
  /* helpers.vhdl:266:50  */
  assign n21411_o = ~n21410_o;
  /* helpers.vhdl:266:46  */
  assign n21412_o = n21409_o & n21411_o;
  /* helpers.vhdl:266:24  */
  assign n21413_o = n21408_o | n21412_o;
  /* helpers.vhdl:266:29  */
  assign n21414_o = n21136_o[39];
  /* helpers.vhdl:266:55  */
  assign n21415_o = n21136_o[35];
  /* helpers.vhdl:266:50  */
  assign n21416_o = ~n21415_o;
  /* helpers.vhdl:266:46  */
  assign n21417_o = n21414_o & n21416_o;
  /* helpers.vhdl:266:24  */
  assign n21418_o = n21413_o | n21417_o;
  /* helpers.vhdl:266:29  */
  assign n21419_o = n21136_o[47];
  /* helpers.vhdl:266:55  */
  assign n21420_o = n21136_o[43];
  /* helpers.vhdl:266:50  */
  assign n21421_o = ~n21420_o;
  /* helpers.vhdl:266:46  */
  assign n21422_o = n21419_o & n21421_o;
  /* helpers.vhdl:266:24  */
  assign n21423_o = n21418_o | n21422_o;
  /* helpers.vhdl:266:29  */
  assign n21424_o = n21136_o[55];
  /* helpers.vhdl:266:55  */
  assign n21425_o = n21136_o[51];
  /* helpers.vhdl:266:50  */
  assign n21426_o = ~n21425_o;
  /* helpers.vhdl:266:46  */
  assign n21427_o = n21424_o & n21426_o;
  /* helpers.vhdl:266:24  */
  assign n21428_o = n21423_o | n21427_o;
  /* helpers.vhdl:266:29  */
  assign n21429_o = n21136_o[63];
  /* helpers.vhdl:266:55  */
  assign n21430_o = n21136_o[59];
  /* helpers.vhdl:266:50  */
  assign n21431_o = ~n21430_o;
  /* helpers.vhdl:266:46  */
  assign n21432_o = n21429_o & n21431_o;
  /* helpers.vhdl:266:24  */
  assign n21433_o = n21428_o | n21432_o;
  /* helpers.vhdl:266:29  */
  assign n21435_o = n21136_o[15];
  /* helpers.vhdl:266:55  */
  assign n21436_o = n21136_o[7];
  /* helpers.vhdl:266:50  */
  assign n21437_o = ~n21436_o;
  /* helpers.vhdl:266:46  */
  assign n21438_o = n21435_o & n21437_o;
  /* helpers.vhdl:266:24  */
  assign n21440_o = 1'b0 | n21438_o;
  /* helpers.vhdl:266:29  */
  assign n21442_o = n21136_o[31];
  /* helpers.vhdl:266:55  */
  assign n21443_o = n21136_o[23];
  /* helpers.vhdl:266:50  */
  assign n21444_o = ~n21443_o;
  /* helpers.vhdl:266:46  */
  assign n21445_o = n21442_o & n21444_o;
  /* helpers.vhdl:266:24  */
  assign n21446_o = n21440_o | n21445_o;
  /* helpers.vhdl:266:29  */
  assign n21447_o = n21136_o[47];
  /* helpers.vhdl:266:55  */
  assign n21448_o = n21136_o[39];
  /* helpers.vhdl:266:50  */
  assign n21449_o = ~n21448_o;
  /* helpers.vhdl:266:46  */
  assign n21450_o = n21447_o & n21449_o;
  /* helpers.vhdl:266:24  */
  assign n21451_o = n21446_o | n21450_o;
  /* helpers.vhdl:266:29  */
  assign n21452_o = n21136_o[63];
  /* helpers.vhdl:266:55  */
  assign n21453_o = n21136_o[55];
  /* helpers.vhdl:266:50  */
  assign n21454_o = ~n21453_o;
  /* helpers.vhdl:266:46  */
  assign n21455_o = n21452_o & n21454_o;
  /* helpers.vhdl:266:24  */
  assign n21456_o = n21451_o | n21455_o;
  /* helpers.vhdl:266:29  */
  assign n21458_o = n21136_o[31];
  /* helpers.vhdl:266:55  */
  assign n21459_o = n21136_o[15];
  /* helpers.vhdl:266:50  */
  assign n21460_o = ~n21459_o;
  /* helpers.vhdl:266:46  */
  assign n21461_o = n21458_o & n21460_o;
  /* helpers.vhdl:266:24  */
  assign n21463_o = 1'b0 | n21461_o;
  /* helpers.vhdl:266:29  */
  assign n21465_o = n21136_o[63];
  /* helpers.vhdl:266:55  */
  assign n21466_o = n21136_o[47];
  /* helpers.vhdl:266:50  */
  assign n21467_o = ~n21466_o;
  /* helpers.vhdl:266:46  */
  assign n21468_o = n21465_o & n21467_o;
  /* helpers.vhdl:266:24  */
  assign n21469_o = n21463_o | n21468_o;
  /* helpers.vhdl:266:29  */
  assign n21471_o = n21136_o[63];
  /* helpers.vhdl:266:55  */
  assign n21472_o = n21136_o[31];
  /* helpers.vhdl:266:50  */
  assign n21473_o = ~n21472_o;
  /* helpers.vhdl:266:46  */
  assign n21474_o = n21471_o & n21473_o;
  /* helpers.vhdl:266:24  */
  assign n21476_o = 1'b0 | n21474_o;
  assign n21478_o = {n21476_o, n21469_o, n21456_o, n21433_o, n21390_o, n21306_o};
  /* helpers.vhdl:286:46  */
  assign n21481_o = {41'b0, n21131_o};  //  uext
  /* helpers.vhdl:244:36  */
  assign n21490_o = n21481_o[1];
  /* helpers.vhdl:244:32  */
  assign n21491_o = |(n21490_o);
  /* helpers.vhdl:244:28  */
  assign n21493_o = 1'b0 | n21491_o;
  /* helpers.vhdl:244:36  */
  assign n21495_o = n21481_o[3];
  /* helpers.vhdl:244:32  */
  assign n21496_o = |(n21495_o);
  /* helpers.vhdl:244:28  */
  assign n21497_o = n21493_o | n21496_o;
  /* helpers.vhdl:244:36  */
  assign n21498_o = n21481_o[5];
  /* helpers.vhdl:244:32  */
  assign n21499_o = |(n21498_o);
  /* helpers.vhdl:244:28  */
  assign n21500_o = n21497_o | n21499_o;
  /* helpers.vhdl:244:36  */
  assign n21501_o = n21481_o[7];
  /* helpers.vhdl:244:32  */
  assign n21502_o = |(n21501_o);
  /* helpers.vhdl:244:28  */
  assign n21503_o = n21500_o | n21502_o;
  /* helpers.vhdl:244:36  */
  assign n21504_o = n21481_o[9];
  /* helpers.vhdl:244:32  */
  assign n21505_o = |(n21504_o);
  /* helpers.vhdl:244:28  */
  assign n21506_o = n21503_o | n21505_o;
  /* helpers.vhdl:244:36  */
  assign n21507_o = n21481_o[11];
  /* helpers.vhdl:244:32  */
  assign n21508_o = |(n21507_o);
  /* helpers.vhdl:244:28  */
  assign n21509_o = n21506_o | n21508_o;
  /* helpers.vhdl:244:36  */
  assign n21510_o = n21481_o[13];
  /* helpers.vhdl:244:32  */
  assign n21511_o = |(n21510_o);
  /* helpers.vhdl:244:28  */
  assign n21512_o = n21509_o | n21511_o;
  /* helpers.vhdl:244:36  */
  assign n21513_o = n21481_o[15];
  /* helpers.vhdl:244:32  */
  assign n21514_o = |(n21513_o);
  /* helpers.vhdl:244:28  */
  assign n21515_o = n21512_o | n21514_o;
  /* helpers.vhdl:244:36  */
  assign n21516_o = n21481_o[17];
  /* helpers.vhdl:244:32  */
  assign n21517_o = |(n21516_o);
  /* helpers.vhdl:244:28  */
  assign n21518_o = n21515_o | n21517_o;
  /* helpers.vhdl:244:36  */
  assign n21519_o = n21481_o[19];
  /* helpers.vhdl:244:32  */
  assign n21520_o = |(n21519_o);
  /* helpers.vhdl:244:28  */
  assign n21521_o = n21518_o | n21520_o;
  /* helpers.vhdl:244:36  */
  assign n21522_o = n21481_o[21];
  /* helpers.vhdl:244:32  */
  assign n21523_o = |(n21522_o);
  /* helpers.vhdl:244:28  */
  assign n21524_o = n21521_o | n21523_o;
  /* helpers.vhdl:244:36  */
  assign n21525_o = n21481_o[23];
  /* helpers.vhdl:244:32  */
  assign n21526_o = |(n21525_o);
  /* helpers.vhdl:244:28  */
  assign n21527_o = n21524_o | n21526_o;
  /* helpers.vhdl:244:36  */
  assign n21528_o = n21481_o[25];
  /* helpers.vhdl:244:32  */
  assign n21529_o = |(n21528_o);
  /* helpers.vhdl:244:28  */
  assign n21530_o = n21527_o | n21529_o;
  /* helpers.vhdl:244:36  */
  assign n21531_o = n21481_o[27];
  /* helpers.vhdl:244:32  */
  assign n21532_o = |(n21531_o);
  /* helpers.vhdl:244:28  */
  assign n21533_o = n21530_o | n21532_o;
  /* helpers.vhdl:244:36  */
  assign n21534_o = n21481_o[29];
  /* helpers.vhdl:244:32  */
  assign n21535_o = |(n21534_o);
  /* helpers.vhdl:244:28  */
  assign n21536_o = n21533_o | n21535_o;
  /* helpers.vhdl:244:36  */
  assign n21537_o = n21481_o[31];
  /* helpers.vhdl:244:32  */
  assign n21538_o = |(n21537_o);
  /* helpers.vhdl:244:28  */
  assign n21539_o = n21536_o | n21538_o;
  /* helpers.vhdl:244:36  */
  assign n21540_o = n21481_o[33];
  /* helpers.vhdl:244:32  */
  assign n21541_o = |(n21540_o);
  /* helpers.vhdl:244:28  */
  assign n21542_o = n21539_o | n21541_o;
  /* helpers.vhdl:244:36  */
  assign n21543_o = n21481_o[35];
  /* helpers.vhdl:244:32  */
  assign n21544_o = |(n21543_o);
  /* helpers.vhdl:244:28  */
  assign n21545_o = n21542_o | n21544_o;
  /* helpers.vhdl:244:36  */
  assign n21546_o = n21481_o[37];
  /* helpers.vhdl:244:32  */
  assign n21547_o = |(n21546_o);
  /* helpers.vhdl:244:28  */
  assign n21548_o = n21545_o | n21547_o;
  /* helpers.vhdl:244:36  */
  assign n21549_o = n21481_o[39];
  /* helpers.vhdl:244:32  */
  assign n21550_o = |(n21549_o);
  /* helpers.vhdl:244:28  */
  assign n21551_o = n21548_o | n21550_o;
  /* helpers.vhdl:244:36  */
  assign n21552_o = n21481_o[41];
  /* helpers.vhdl:244:32  */
  assign n21553_o = |(n21552_o);
  /* helpers.vhdl:244:28  */
  assign n21554_o = n21551_o | n21553_o;
  /* helpers.vhdl:244:36  */
  assign n21555_o = n21481_o[43];
  /* helpers.vhdl:244:32  */
  assign n21556_o = |(n21555_o);
  /* helpers.vhdl:244:28  */
  assign n21557_o = n21554_o | n21556_o;
  /* helpers.vhdl:244:36  */
  assign n21558_o = n21481_o[45];
  /* helpers.vhdl:244:32  */
  assign n21559_o = |(n21558_o);
  /* helpers.vhdl:244:28  */
  assign n21560_o = n21557_o | n21559_o;
  /* helpers.vhdl:244:36  */
  assign n21561_o = n21481_o[47];
  /* helpers.vhdl:244:32  */
  assign n21562_o = |(n21561_o);
  /* helpers.vhdl:244:28  */
  assign n21563_o = n21560_o | n21562_o;
  /* helpers.vhdl:244:36  */
  assign n21564_o = n21481_o[49];
  /* helpers.vhdl:244:32  */
  assign n21565_o = |(n21564_o);
  /* helpers.vhdl:244:28  */
  assign n21566_o = n21563_o | n21565_o;
  /* helpers.vhdl:244:36  */
  assign n21567_o = n21481_o[51];
  /* helpers.vhdl:244:32  */
  assign n21568_o = |(n21567_o);
  /* helpers.vhdl:244:28  */
  assign n21569_o = n21566_o | n21568_o;
  /* helpers.vhdl:244:36  */
  assign n21570_o = n21481_o[53];
  /* helpers.vhdl:244:32  */
  assign n21571_o = |(n21570_o);
  /* helpers.vhdl:244:28  */
  assign n21572_o = n21569_o | n21571_o;
  /* helpers.vhdl:244:36  */
  assign n21573_o = n21481_o[55];
  /* helpers.vhdl:244:32  */
  assign n21574_o = |(n21573_o);
  /* helpers.vhdl:244:28  */
  assign n21575_o = n21572_o | n21574_o;
  /* helpers.vhdl:244:36  */
  assign n21576_o = n21481_o[57];
  /* helpers.vhdl:244:32  */
  assign n21577_o = |(n21576_o);
  /* helpers.vhdl:244:28  */
  assign n21578_o = n21575_o | n21577_o;
  /* helpers.vhdl:244:36  */
  assign n21579_o = n21481_o[59];
  /* helpers.vhdl:244:32  */
  assign n21580_o = |(n21579_o);
  /* helpers.vhdl:244:28  */
  assign n21581_o = n21578_o | n21580_o;
  /* helpers.vhdl:244:36  */
  assign n21582_o = n21481_o[61];
  /* helpers.vhdl:244:32  */
  assign n21583_o = |(n21582_o);
  /* helpers.vhdl:244:28  */
  assign n21584_o = n21581_o | n21583_o;
  /* helpers.vhdl:244:36  */
  assign n21585_o = n21481_o[63];
  /* helpers.vhdl:244:32  */
  assign n21586_o = |(n21585_o);
  /* helpers.vhdl:244:28  */
  assign n21587_o = n21584_o | n21586_o;
  /* helpers.vhdl:244:36  */
  assign n21590_o = n21481_o[3:2];
  /* helpers.vhdl:244:32  */
  assign n21591_o = |(n21590_o);
  /* helpers.vhdl:244:28  */
  assign n21593_o = 1'b0 | n21591_o;
  /* helpers.vhdl:244:36  */
  assign n21595_o = n21481_o[7:6];
  /* helpers.vhdl:244:32  */
  assign n21596_o = |(n21595_o);
  /* helpers.vhdl:244:28  */
  assign n21597_o = n21593_o | n21596_o;
  /* helpers.vhdl:244:36  */
  assign n21598_o = n21481_o[11:10];
  /* helpers.vhdl:244:32  */
  assign n21599_o = |(n21598_o);
  /* helpers.vhdl:244:28  */
  assign n21600_o = n21597_o | n21599_o;
  /* helpers.vhdl:244:36  */
  assign n21601_o = n21481_o[15:14];
  /* helpers.vhdl:244:32  */
  assign n21602_o = |(n21601_o);
  /* helpers.vhdl:244:28  */
  assign n21603_o = n21600_o | n21602_o;
  /* helpers.vhdl:244:36  */
  assign n21604_o = n21481_o[19:18];
  /* helpers.vhdl:244:32  */
  assign n21605_o = |(n21604_o);
  /* helpers.vhdl:244:28  */
  assign n21606_o = n21603_o | n21605_o;
  /* helpers.vhdl:244:36  */
  assign n21607_o = n21481_o[23:22];
  /* helpers.vhdl:244:32  */
  assign n21608_o = |(n21607_o);
  /* helpers.vhdl:244:28  */
  assign n21609_o = n21606_o | n21608_o;
  /* helpers.vhdl:244:36  */
  assign n21610_o = n21481_o[27:26];
  /* helpers.vhdl:244:32  */
  assign n21611_o = |(n21610_o);
  /* helpers.vhdl:244:28  */
  assign n21612_o = n21609_o | n21611_o;
  /* helpers.vhdl:244:36  */
  assign n21613_o = n21481_o[31:30];
  /* helpers.vhdl:244:32  */
  assign n21614_o = |(n21613_o);
  /* helpers.vhdl:244:28  */
  assign n21615_o = n21612_o | n21614_o;
  /* helpers.vhdl:244:36  */
  assign n21616_o = n21481_o[35:34];
  /* helpers.vhdl:244:32  */
  assign n21617_o = |(n21616_o);
  /* helpers.vhdl:244:28  */
  assign n21618_o = n21615_o | n21617_o;
  /* helpers.vhdl:244:36  */
  assign n21619_o = n21481_o[39:38];
  /* helpers.vhdl:244:32  */
  assign n21620_o = |(n21619_o);
  /* helpers.vhdl:244:28  */
  assign n21621_o = n21618_o | n21620_o;
  /* helpers.vhdl:244:36  */
  assign n21622_o = n21481_o[43:42];
  /* helpers.vhdl:244:32  */
  assign n21623_o = |(n21622_o);
  /* helpers.vhdl:244:28  */
  assign n21624_o = n21621_o | n21623_o;
  /* helpers.vhdl:244:36  */
  assign n21625_o = n21481_o[47:46];
  /* helpers.vhdl:244:32  */
  assign n21626_o = |(n21625_o);
  /* helpers.vhdl:244:28  */
  assign n21627_o = n21624_o | n21626_o;
  /* helpers.vhdl:244:36  */
  assign n21628_o = n21481_o[51:50];
  /* helpers.vhdl:244:32  */
  assign n21629_o = |(n21628_o);
  /* helpers.vhdl:244:28  */
  assign n21630_o = n21627_o | n21629_o;
  /* helpers.vhdl:244:36  */
  assign n21631_o = n21481_o[55:54];
  /* helpers.vhdl:244:32  */
  assign n21632_o = |(n21631_o);
  /* helpers.vhdl:244:28  */
  assign n21633_o = n21630_o | n21632_o;
  /* helpers.vhdl:244:36  */
  assign n21634_o = n21481_o[59:58];
  /* helpers.vhdl:244:32  */
  assign n21635_o = |(n21634_o);
  /* helpers.vhdl:244:28  */
  assign n21636_o = n21633_o | n21635_o;
  /* helpers.vhdl:244:36  */
  assign n21637_o = n21481_o[63:62];
  /* helpers.vhdl:244:32  */
  assign n21638_o = |(n21637_o);
  /* helpers.vhdl:244:28  */
  assign n21639_o = n21636_o | n21638_o;
  /* helpers.vhdl:244:36  */
  assign n21641_o = n21481_o[7:4];
  /* helpers.vhdl:244:32  */
  assign n21642_o = |(n21641_o);
  /* helpers.vhdl:244:28  */
  assign n21644_o = 1'b0 | n21642_o;
  /* helpers.vhdl:244:36  */
  assign n21646_o = n21481_o[15:12];
  /* helpers.vhdl:244:32  */
  assign n21647_o = |(n21646_o);
  /* helpers.vhdl:244:28  */
  assign n21648_o = n21644_o | n21647_o;
  /* helpers.vhdl:244:36  */
  assign n21649_o = n21481_o[23:20];
  /* helpers.vhdl:244:32  */
  assign n21650_o = |(n21649_o);
  /* helpers.vhdl:244:28  */
  assign n21651_o = n21648_o | n21650_o;
  /* helpers.vhdl:244:36  */
  assign n21652_o = n21481_o[31:28];
  /* helpers.vhdl:244:32  */
  assign n21653_o = |(n21652_o);
  /* helpers.vhdl:244:28  */
  assign n21654_o = n21651_o | n21653_o;
  /* helpers.vhdl:244:36  */
  assign n21655_o = n21481_o[39:36];
  /* helpers.vhdl:244:32  */
  assign n21656_o = |(n21655_o);
  /* helpers.vhdl:244:28  */
  assign n21657_o = n21654_o | n21656_o;
  /* helpers.vhdl:244:36  */
  assign n21658_o = n21481_o[47:44];
  /* helpers.vhdl:244:32  */
  assign n21659_o = |(n21658_o);
  /* helpers.vhdl:244:28  */
  assign n21660_o = n21657_o | n21659_o;
  /* helpers.vhdl:244:36  */
  assign n21661_o = n21481_o[55:52];
  /* helpers.vhdl:244:32  */
  assign n21662_o = |(n21661_o);
  /* helpers.vhdl:244:28  */
  assign n21663_o = n21660_o | n21662_o;
  /* helpers.vhdl:244:36  */
  assign n21664_o = n21481_o[63:60];
  /* helpers.vhdl:244:32  */
  assign n21665_o = |(n21664_o);
  /* helpers.vhdl:244:28  */
  assign n21666_o = n21663_o | n21665_o;
  /* helpers.vhdl:244:36  */
  assign n21668_o = n21481_o[15:8];
  /* helpers.vhdl:244:32  */
  assign n21669_o = |(n21668_o);
  /* helpers.vhdl:244:28  */
  assign n21671_o = 1'b0 | n21669_o;
  /* helpers.vhdl:244:36  */
  assign n21673_o = n21481_o[31:24];
  /* helpers.vhdl:244:32  */
  assign n21674_o = |(n21673_o);
  /* helpers.vhdl:244:28  */
  assign n21675_o = n21671_o | n21674_o;
  /* helpers.vhdl:244:36  */
  assign n21676_o = n21481_o[47:40];
  /* helpers.vhdl:244:32  */
  assign n21677_o = |(n21676_o);
  /* helpers.vhdl:244:28  */
  assign n21678_o = n21675_o | n21677_o;
  /* helpers.vhdl:244:36  */
  assign n21679_o = n21481_o[63:56];
  /* helpers.vhdl:244:32  */
  assign n21680_o = |(n21679_o);
  /* helpers.vhdl:244:28  */
  assign n21681_o = n21678_o | n21680_o;
  /* helpers.vhdl:244:36  */
  assign n21683_o = n21481_o[31:16];
  /* helpers.vhdl:244:32  */
  assign n21684_o = |(n21683_o);
  /* helpers.vhdl:244:28  */
  assign n21686_o = 1'b0 | n21684_o;
  /* helpers.vhdl:244:36  */
  assign n21688_o = n21481_o[63:48];
  /* helpers.vhdl:244:32  */
  assign n21689_o = |(n21688_o);
  /* helpers.vhdl:244:28  */
  assign n21690_o = n21686_o | n21689_o;
  /* helpers.vhdl:244:36  */
  assign n21692_o = n21481_o[63:32];
  /* helpers.vhdl:244:32  */
  assign n21693_o = |(n21692_o);
  /* helpers.vhdl:244:28  */
  assign n21695_o = 1'b0 | n21693_o;
  assign n21697_o = {n21695_o, n21690_o, n21681_o, n21666_o, n21639_o, n21587_o};
  /* helpers.vhdl:287:19  */
  assign n21699_o = n21478_o[5:2];
  /* helpers.vhdl:287:38  */
  assign n21700_o = n21697_o[1:0];
  /* helpers.vhdl:287:32  */
  assign n21701_o = {n21699_o, n21700_o};
  /* loadstore1.vhdl:735:17  */
  assign n21704_o = n19358_o[0];
  /* loadstore1.vhdl:735:36  */
  assign n21705_o = r2[272:0];
  /* loadstore1.vhdl:735:40  */
  assign n21706_o = n21705_o[2];
  /* loadstore1.vhdl:735:29  */
  assign n21707_o = n21704_o & n21706_o;
  assign n21708_o = {n22420_o, n22406_o, n22392_o, n22378_o, n22364_o, n22350_o, n22336_o, n22322_o};
  assign n21709_o = r3[148:85];
  /* loadstore1.vhdl:735:9  */
  assign n21710_o = n21707_o ? n21708_o : n21709_o;
  assign n21711_o = r3[244:149];
  /* loadstore1.vhdl:739:15  */
  assign n21712_o = r2[272:0];
  /* loadstore1.vhdl:739:19  */
  assign n21713_o = n21712_o[0];
  /* loadstore1.vhdl:740:19  */
  assign n21714_o = r2[272:0];
  /* loadstore1.vhdl:740:23  */
  assign n21715_o = n21714_o[6];
  /* loadstore1.vhdl:744:31  */
  assign n21716_o = r2[203];
  /* loadstore1.vhdl:744:35  */
  assign n21717_o = ~n21716_o;
  /* loadstore1.vhdl:744:56  */
  assign n21718_o = r2[200];
  /* loadstore1.vhdl:744:60  */
  assign n21719_o = ~n21718_o;
  /* loadstore1.vhdl:744:41  */
  assign n21720_o = n21717_o & n21719_o;
  /* loadstore1.vhdl:745:35  */
  assign n21721_o = r2[195];
  /* loadstore1.vhdl:745:39  */
  assign n21722_o = ~n21721_o;
  /* loadstore1.vhdl:746:52  */
  assign n21723_o = r3[244:213];
  /* loadstore1.vhdl:746:47  */
  assign n21725_o = {32'b00000000000000000000000000000000, n21723_o};
  /* loadstore1.vhdl:748:38  */
  assign n21726_o = r3[212:149];
  /* loadstore1.vhdl:745:21  */
  assign n21727_o = n21722_o ? n21725_o : n21726_o;
  /* loadstore1.vhdl:752:36  */
  assign n21728_o = n19370_o[70:7];
  /* loadstore1.vhdl:744:17  */
  assign n21729_o = n21720_o ? n21727_o : n21728_o;
  /* loadstore1.vhdl:740:13  */
  assign n21732_o = n21715_o ? 1'b1 : 1'b0;
  /* loadstore1.vhdl:740:13  */
  assign n21734_o = n21715_o ? n21729_o : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* loadstore1.vhdl:755:19  */
  assign n21735_o = r2[272:0];
  /* loadstore1.vhdl:755:23  */
  assign n21736_o = n21735_o[206];
  /* loadstore1.vhdl:755:13  */
  assign n21739_o = n21736_o ? 1'b1 : 1'b0;
  /* loadstore1.vhdl:759:19  */
  assign n21740_o = r2[272:0];
  /* loadstore1.vhdl:759:23  */
  assign n21741_o = n21740_o[10];
  /* loadstore1.vhdl:759:13  */
  assign n21743_o = n21741_o ? 1'b1 : n21732_o;
  /* loadstore1.vhdl:762:19  */
  assign n21744_o = r2[272:0];
  /* loadstore1.vhdl:762:23  */
  assign n21745_o = n21744_o[11];
  /* loadstore1.vhdl:762:13  */
  assign n21748_o = n21745_o ? 1'b1 : 1'b0;
  /* loadstore1.vhdl:739:9  */
  assign n21750_o = n21713_o ? n21743_o : 1'b0;
  /* loadstore1.vhdl:739:9  */
  assign n21753_o = n21713_o ? n21748_o : 1'b0;
  /* loadstore1.vhdl:739:9  */
  assign n21756_o = n21713_o ? n21739_o : 1'b0;
  /* loadstore1.vhdl:739:9  */
  assign n21759_o = n21713_o ? n21734_o : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* loadstore1.vhdl:767:17  */
  assign n21761_o = r3[1:0];
  /* loadstore1.vhdl:769:21  */
  assign n21762_o = n19358_o[0];
  /* loadstore1.vhdl:770:23  */
  assign n21763_o = r2[272:0];
  /* loadstore1.vhdl:770:27  */
  assign n21764_o = n21763_o[208];
  /* loadstore1.vhdl:770:38  */
  assign n21765_o = ~n21764_o;
  /* loadstore1.vhdl:770:50  */
  assign n21766_o = r2[272:0];
  /* loadstore1.vhdl:770:54  */
  assign n21767_o = n21766_o[207];
  /* loadstore1.vhdl:770:44  */
  assign n21768_o = n21765_o | n21767_o;
  /* loadstore1.vhdl:771:40  */
  assign n21769_o = r2[272:0];
  /* loadstore1.vhdl:771:44  */
  assign n21770_o = n21769_o[2];
  /* loadstore1.vhdl:771:60  */
  assign n21771_o = r2[272:0];
  /* loadstore1.vhdl:771:64  */
  assign n21772_o = n21771_o[194];
  /* loadstore1.vhdl:771:53  */
  assign n21773_o = ~n21772_o;
  /* loadstore1.vhdl:771:49  */
  assign n21774_o = n21770_o & n21773_o;
  /* loadstore1.vhdl:772:39  */
  assign n21775_o = r2[272:0];
  /* loadstore1.vhdl:772:43  */
  assign n21776_o = n21775_o[194];
  /* loadstore1.vhdl:772:32  */
  assign n21778_o = 1'b1 & n21776_o;
  /* loadstore1.vhdl:778:41  */
  assign n21781_o = r2[272:0];
  /* loadstore1.vhdl:778:45  */
  assign n21782_o = n21781_o[181];
  /* loadstore1.vhdl:778:59  */
  assign n21783_o = r2[272:0];
  /* loadstore1.vhdl:778:63  */
  assign n21784_o = n21783_o[3];
  /* loadstore1.vhdl:778:52  */
  assign n21785_o = n21782_o & n21784_o;
  assign n21786_o = r3[1:0];
  /* loadstore1.vhdl:769:13  */
  assign n21787_o = n21799_o ? 2'b11 : n21786_o;
  /* loadstore1.vhdl:769:13  */
  assign n21788_o = n21800_o ? 1'b1 : 1'b0;
  /* loadstore1.vhdl:772:21  */
  assign n21789_o = n21778_o ? n21753_o : n21785_o;
  /* loadstore1.vhdl:770:17  */
  assign n21791_o = n21768_o & n21778_o;
  /* loadstore1.vhdl:770:17  */
  assign n21792_o = n21768_o & n21778_o;
  /* loadstore1.vhdl:769:13  */
  assign n21793_o = n21801_o ? n21774_o : n21750_o;
  /* loadstore1.vhdl:769:13  */
  assign n21794_o = n21802_o ? n21789_o : n21753_o;
  /* loadstore1.vhdl:770:17  */
  assign n21797_o = n21768_o ? 1'b0 : 1'b1;
  /* loadstore1.vhdl:769:13  */
  assign n21799_o = n21762_o & n21791_o;
  /* loadstore1.vhdl:769:13  */
  assign n21800_o = n21762_o & n21792_o;
  /* loadstore1.vhdl:769:13  */
  assign n21801_o = n21762_o & n21768_o;
  /* loadstore1.vhdl:769:13  */
  assign n21802_o = n21762_o & n21768_o;
  /* loadstore1.vhdl:769:13  */
  assign n21804_o = n21762_o ? n21797_o : 1'b0;
  /* loadstore1.vhdl:784:21  */
  assign n21805_o = n19358_o[66];
  /* loadstore1.vhdl:785:25  */
  assign n21806_o = n19358_o[67];
  /* loadstore1.vhdl:788:46  */
  assign n21807_o = r2[272:0];
  /* loadstore1.vhdl:788:50  */
  assign n21808_o = n21807_o[2];
  /* loadstore1.vhdl:788:39  */
  assign n21809_o = ~n21808_o;
  /* loadstore1.vhdl:791:44  */
  assign n21810_o = n19358_o[67];
  /* loadstore1.vhdl:785:17  */
  assign n21813_o = n21806_o ? n21787_o : 2'b01;
  assign n21814_o = r3[284];
  /* loadstore1.vhdl:785:17  */
  assign n21815_o = n21806_o ? n21814_o : 1'b0;
  /* loadstore1.vhdl:785:17  */
  assign n21818_o = n21806_o ? 1'b0 : 1'b1;
  /* loadstore1.vhdl:784:13  */
  assign n21820_o = n21830_o ? 1'b1 : n21756_o;
  /* loadstore1.vhdl:785:17  */
  assign n21822_o = n21806_o ? n21809_o : 1'b0;
  /* loadstore1.vhdl:785:17  */
  assign n21824_o = n21806_o ? n21810_o : 1'b0;
  /* loadstore1.vhdl:784:13  */
  assign n21825_o = n21805_o ? n21813_o : n21787_o;
  assign n21826_o = r3[284];
  /* loadstore1.vhdl:784:13  */
  assign n21827_o = n21805_o ? n21815_o : n21826_o;
  /* loadstore1.vhdl:784:13  */
  assign n21829_o = n21805_o ? n21818_o : 1'b0;
  /* loadstore1.vhdl:784:13  */
  assign n21830_o = n21805_o & n21806_o;
  /* loadstore1.vhdl:784:13  */
  assign n21832_o = n21805_o ? n21822_o : 1'b0;
  /* loadstore1.vhdl:784:13  */
  assign n21834_o = n21805_o ? n21824_o : 1'b0;
  /* loadstore1.vhdl:801:19  */
  assign n21835_o = r2[272:0];
  /* loadstore1.vhdl:801:23  */
  assign n21836_o = n21835_o[0];
  /* loadstore1.vhdl:802:23  */
  assign n21837_o = r2[272:0];
  /* loadstore1.vhdl:802:27  */
  assign n21838_o = n21837_o[8];
  /* loadstore1.vhdl:804:38  */
  assign n21839_o = r2[272:0];
  /* loadstore1.vhdl:804:42  */
  assign n21840_o = n21839_o[7];
  /* loadstore1.vhdl:804:31  */
  assign n21841_o = ~n21840_o;
  /* loadstore1.vhdl:805:37  */
  assign n21842_o = r2[272:0];
  /* loadstore1.vhdl:805:41  */
  assign n21843_o = n21842_o[7];
  /* loadstore1.vhdl:806:27  */
  assign n21844_o = r2[272:0];
  /* loadstore1.vhdl:806:31  */
  assign n21845_o = n21844_o[9];
  /* loadstore1.vhdl:806:21  */
  assign n21849_o = n21845_o ? 2'b01 : 2'b10;
  assign n21850_o = n20503_o[2];
  /* loadstore1.vhdl:801:13  */
  assign n21851_o = n21875_o ? 1'b1 : n21850_o;
  /* loadstore1.vhdl:812:26  */
  assign n21852_o = r2[272:0];
  /* loadstore1.vhdl:812:30  */
  assign n21853_o = n21852_o[7];
  /* loadstore1.vhdl:813:35  */
  assign n21854_o = r2[195];
  /* loadstore1.vhdl:813:39  */
  assign n21855_o = ~n21854_o;
  /* loadstore1.vhdl:814:53  */
  assign n21856_o = r2[125:94];
  /* loadstore1.vhdl:816:37  */
  assign n21857_o = r2[272:0];
  /* loadstore1.vhdl:816:41  */
  assign n21858_o = n21857_o[157:94];
  assign n21859_o = r3[212:149];
  /* loadstore1.vhdl:813:21  */
  assign n21860_o = n21855_o ? n21859_o : n21858_o;
  assign n21861_o = r3[244:213];
  /* loadstore1.vhdl:813:21  */
  assign n21862_o = n21855_o ? n21856_o : n21861_o;
  assign n21863_o = {n21862_o, n21860_o};
  /* loadstore1.vhdl:812:17  */
  assign n21864_o = n21853_o ? n21863_o : n21711_o;
  /* loadstore1.vhdl:801:13  */
  assign n21865_o = n21872_o ? n21849_o : n21825_o;
  /* loadstore1.vhdl:802:17  */
  assign n21866_o = n21838_o ? n21711_o : n21864_o;
  /* loadstore1.vhdl:802:17  */
  assign n21868_o = n21838_o & n21845_o;
  /* loadstore1.vhdl:801:13  */
  assign n21869_o = n21876_o ? n21841_o : n21829_o;
  /* loadstore1.vhdl:802:17  */
  assign n21871_o = n21838_o ? n21843_o : 1'b0;
  /* loadstore1.vhdl:801:13  */
  assign n21872_o = n21836_o & n21838_o;
  /* loadstore1.vhdl:801:13  */
  assign n21873_o = n21836_o ? n21866_o : n21711_o;
  /* loadstore1.vhdl:801:13  */
  assign n21875_o = n21836_o & n21868_o;
  /* loadstore1.vhdl:801:13  */
  assign n21876_o = n21836_o & n21838_o;
  /* loadstore1.vhdl:801:13  */
  assign n21878_o = n21836_o ? n21871_o : 1'b0;
  /* loadstore1.vhdl:768:9  */
  assign n21880_o = n21761_o == 2'b00;
  /* loadstore1.vhdl:822:21  */
  assign n21881_o = n19370_o[0];
  /* loadstore1.vhdl:823:23  */
  assign n21882_o = r2[272:0];
  /* loadstore1.vhdl:823:27  */
  assign n21883_o = n21882_o[9];
  /* loadstore1.vhdl:823:39  */
  assign n21884_o = ~n21883_o;
  assign n21887_o = r3[1:0];
  /* loadstore1.vhdl:822:13  */
  assign n21888_o = n21895_o ? 2'b00 : n21887_o;
  assign n21889_o = r3[284];
  /* loadstore1.vhdl:822:13  */
  assign n21890_o = n21897_o ? 1'b1 : n21889_o;
  /* loadstore1.vhdl:823:17  */
  assign n21893_o = n21884_o ? 1'b1 : 1'b0;
  /* loadstore1.vhdl:822:13  */
  assign n21895_o = n21881_o & n21884_o;
  /* loadstore1.vhdl:822:13  */
  assign n21897_o = n21881_o & n21884_o;
  /* loadstore1.vhdl:822:13  */
  assign n21899_o = n21881_o ? n21893_o : 1'b0;
  /* loadstore1.vhdl:830:21  */
  assign n21900_o = n19370_o[1];
  /* loadstore1.vhdl:832:40  */
  assign n21901_o = n19370_o[2];
  /* loadstore1.vhdl:833:40  */
  assign n21902_o = n19370_o[5];
  /* loadstore1.vhdl:834:38  */
  assign n21903_o = r2[272:0];
  /* loadstore1.vhdl:834:42  */
  assign n21904_o = n21903_o[3];
  /* loadstore1.vhdl:834:54  */
  assign n21905_o = r2[272:0];
  /* loadstore1.vhdl:834:58  */
  assign n21906_o = n21905_o[5];
  /* loadstore1.vhdl:834:48  */
  assign n21907_o = n21904_o | n21906_o;
  /* loadstore1.vhdl:835:40  */
  assign n21908_o = n19370_o[3];
  /* loadstore1.vhdl:836:40  */
  assign n21909_o = n19370_o[6];
  /* loadstore1.vhdl:830:13  */
  assign n21911_o = n21900_o ? 1'b1 : n21756_o;
  assign n21912_o = {n21908_o, n21909_o};
  /* loadstore1.vhdl:830:13  */
  assign n21914_o = n21900_o ? n21912_o : 2'b00;
  /* loadstore1.vhdl:830:13  */
  assign n21916_o = n21900_o ? n21907_o : 1'b0;
  /* loadstore1.vhdl:830:13  */
  assign n21918_o = n21900_o ? n21902_o : 1'b0;
  /* loadstore1.vhdl:830:13  */
  assign n21920_o = n21900_o ? n21901_o : 1'b0;
  /* loadstore1.vhdl:821:9  */
  assign n21922_o = n21761_o == 2'b01;
  /* loadstore1.vhdl:839:9  */
  assign n21924_o = n21761_o == 2'b10;
  /* loadstore1.vhdl:841:9  */
  assign n21926_o = n21761_o == 2'b11;
  assign n21927_o = {n21926_o, n21924_o, n21922_o, n21880_o};
  assign n21928_o = r3[1:0];
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21930_o = n21928_o;
      4'b0100: n21930_o = n21928_o;
      4'b0010: n21930_o = n21888_o;
      4'b0001: n21930_o = n21865_o;
      default: n21930_o = 2'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21932_o = 1'b0;
      4'b0100: n21932_o = 1'b0;
      4'b0010: n21932_o = 1'b0;
      4'b0001: n21932_o = n21788_o;
      default: n21932_o = 1'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21934_o = n21711_o;
      4'b0100: n21934_o = n21711_o;
      4'b0010: n21934_o = n21711_o;
      4'b0001: n21934_o = n21873_o;
      default: n21934_o = 96'bX;
    endcase
  assign n21935_o = r3[284];
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21937_o = n21935_o;
      4'b0100: n21937_o = n21935_o;
      4'b0010: n21937_o = n21890_o;
      4'b0001: n21937_o = n21827_o;
      default: n21937_o = 1'bX;
    endcase
  assign n21938_o = n20503_o[2];
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21940_o = n21938_o;
      4'b0100: n21940_o = n21938_o;
      4'b0010: n21940_o = n21938_o;
      4'b0001: n21940_o = n21851_o;
      default: n21940_o = 1'bX;
    endcase
  assign n21941_o = r3[83:2];
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21946_o = 1'b0;
      4'b0100: n21946_o = 1'b0;
      4'b0010: n21946_o = n21899_o;
      4'b0001: n21946_o = 1'b0;
      default: n21946_o = 1'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21950_o = 1'b0;
      4'b0100: n21950_o = 1'b0;
      4'b0010: n21950_o = 1'b0;
      4'b0001: n21950_o = n21869_o;
      default: n21950_o = 1'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21954_o = 1'b0;
      4'b0100: n21954_o = 1'b0;
      4'b0010: n21954_o = 1'b0;
      4'b0001: n21954_o = n21878_o;
      default: n21954_o = 1'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21958_o = 1'b1;
      4'b0100: n21958_o = n21750_o;
      4'b0010: n21958_o = n21750_o;
      4'b0001: n21958_o = n21793_o;
      default: n21958_o = 1'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21960_o = n21753_o;
      4'b0100: n21960_o = n21753_o;
      4'b0010: n21960_o = n21753_o;
      4'b0001: n21960_o = n21794_o;
      default: n21960_o = 1'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21963_o = 1'b0;
      4'b0100: n21963_o = 1'b0;
      4'b0010: n21963_o = 1'b0;
      4'b0001: n21963_o = n21804_o;
      default: n21963_o = 1'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21966_o = n21756_o;
      4'b0100: n21966_o = n21756_o;
      4'b0010: n21966_o = n21911_o;
      4'b0001: n21966_o = n21820_o;
      default: n21966_o = 1'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21969_o = 2'b00;
      4'b0100: n21969_o = 2'b00;
      4'b0010: n21969_o = n21914_o;
      4'b0001: n21969_o = 2'b00;
      default: n21969_o = 2'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21972_o = 1'b0;
      4'b0100: n21972_o = 1'b0;
      4'b0010: n21972_o = n21916_o;
      4'b0001: n21972_o = n21832_o;
      default: n21972_o = 1'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21975_o = 1'b0;
      4'b0100: n21975_o = 1'b0;
      4'b0010: n21975_o = n21918_o;
      4'b0001: n21975_o = 1'b0;
      default: n21975_o = 1'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21978_o = 1'b0;
      4'b0100: n21978_o = 1'b0;
      4'b0010: n21978_o = 1'b0;
      4'b0001: n21978_o = n21834_o;
      default: n21978_o = 1'bX;
    endcase
  /* loadstore1.vhdl:767:9  */
  always @*
    case (n21927_o)
      4'b1000: n21981_o = 1'b0;
      4'b0100: n21981_o = 1'b0;
      4'b0010: n21981_o = n21920_o;
      4'b0001: n21981_o = 1'b0;
      default: n21981_o = 1'bX;
    endcase
  assign n21984_o = n21982_o[17:0];
  assign n21986_o = n21982_o[24:20];
  assign n21988_o = n21982_o[26];
  assign n21990_o = n21982_o[31];
  assign n21991_o = n21982_o[29];
  /* loadstore1.vhdl:846:27  */
  assign n21992_o = complete | n21966_o;
  /* loadstore1.vhdl:846:9  */
  assign n21995_o = n21992_o ? 2'b00 : n21930_o;
  /* loadstore1.vhdl:846:9  */
  assign n21996_o = n21992_o ? 1'b1 : n21937_o;
  /* loadstore1.vhdl:851:38  */
  assign n21997_o = r2[272:0];
  /* loadstore1.vhdl:851:42  */
  assign n21998_o = n21997_o[2];
  /* loadstore1.vhdl:851:47  */
  assign n21999_o = n21998_o & complete;
  /* loadstore1.vhdl:852:40  */
  assign n22001_o = r2[272:0];
  /* loadstore1.vhdl:852:44  */
  assign n22002_o = n22001_o[3];
  /* loadstore1.vhdl:852:56  */
  assign n22003_o = r2[272:0];
  /* loadstore1.vhdl:852:60  */
  assign n22004_o = n22003_o[5];
  /* loadstore1.vhdl:852:50  */
  assign n22005_o = n22002_o | n22004_o;
  /* loadstore1.vhdl:852:66  */
  assign n22006_o = n22005_o & complete;
  assign n22007_o = r3[361:286];
  /* loadstore1.vhdl:858:25  */
  assign n22008_o = r2[272:0];
  /* loadstore1.vhdl:858:29  */
  assign n22009_o = n22008_o[272:209];
  /* loadstore1.vhdl:859:19  */
  assign n22010_o = r2[272:0];
  /* loadstore1.vhdl:859:23  */
  assign n22011_o = n22010_o[206];
  /* loadstore1.vhdl:861:29  */
  assign n22013_o = r2[272:0];
  /* loadstore1.vhdl:861:33  */
  assign n22014_o = n22013_o[77:14];
  /* loadstore1.vhdl:862:22  */
  assign n22015_o = r2[272:0];
  /* loadstore1.vhdl:862:26  */
  assign n22016_o = n22015_o[9];
  /* loadstore1.vhdl:862:38  */
  assign n22017_o = ~n22016_o;
  /* loadstore1.vhdl:863:29  */
  assign n22018_o = r2[272:0];
  /* loadstore1.vhdl:863:33  */
  assign n22019_o = n22018_o[77:14];
  /* loadstore1.vhdl:864:25  */
  assign n22020_o = n19370_o[4];
  /* loadstore1.vhdl:864:32  */
  assign n22021_o = ~n22020_o;
  assign n22023_o = {n21990_o, n21981_o, n21991_o, n21978_o, n21975_o, n21988_o, n21972_o, n21986_o, n21969_o, n21984_o};
  assign n22025_o = n21934_o[95:64];
  /* loadstore1.vhdl:864:17  */
  assign n22026_o = n22021_o ? n22023_o : n22025_o;
  /* loadstore1.vhdl:864:17  */
  assign n22027_o = n22021_o ? 12'b001100000000 : 12'b001110000000;
  /* loadstore1.vhdl:871:25  */
  assign n22028_o = n19370_o[4];
  /* loadstore1.vhdl:871:32  */
  assign n22029_o = ~n22028_o;
  /* loadstore1.vhdl:872:45  */
  assign n22030_o = n19370_o[2];
  /* loadstore1.vhdl:873:45  */
  assign n22031_o = n19370_o[5];
  /* loadstore1.vhdl:874:45  */
  assign n22032_o = n19370_o[3];
  /* loadstore1.vhdl:875:45  */
  assign n22033_o = n19370_o[6];
  assign n22036_o = {n22032_o, n22033_o};
  /* loadstore1.vhdl:871:17  */
  assign n22037_o = n22029_o ? 12'b010000000000 : 12'b010010000000;
  assign n22038_o = n20500_o[3:2];
  /* loadstore1.vhdl:871:17  */
  assign n22039_o = n22029_o ? n22036_o : n22038_o;
  assign n22040_o = n20500_o[12];
  /* loadstore1.vhdl:871:17  */
  assign n22041_o = n22029_o ? n22031_o : n22040_o;
  assign n22042_o = n20500_o[14];
  /* loadstore1.vhdl:871:17  */
  assign n22043_o = n22029_o ? n22030_o : n22042_o;
  assign n22044_o = {n22026_o, n22019_o};
  /* loadstore1.vhdl:862:13  */
  assign n22045_o = n22017_o ? n22044_o : n21934_o;
  /* loadstore1.vhdl:862:13  */
  assign n22046_o = n22017_o ? n22027_o : n22037_o;
  assign n22047_o = n20500_o[3:2];
  /* loadstore1.vhdl:862:13  */
  assign n22048_o = n22017_o ? n22047_o : n22039_o;
  assign n22049_o = n20500_o[12];
  /* loadstore1.vhdl:862:13  */
  assign n22050_o = n22017_o ? n22049_o : n22041_o;
  assign n22051_o = n20500_o[14];
  /* loadstore1.vhdl:862:13  */
  assign n22052_o = n22017_o ? n22051_o : n22043_o;
  assign n22053_o = n22045_o[63:0];
  /* loadstore1.vhdl:859:13  */
  assign n22054_o = n22011_o ? n22014_o : n22053_o;
  assign n22055_o = n22045_o[95:64];
  assign n22056_o = n21934_o[95:64];
  /* loadstore1.vhdl:859:13  */
  assign n22057_o = n22011_o ? n22056_o : n22055_o;
  /* loadstore1.vhdl:859:13  */
  assign n22058_o = n22011_o ? 12'b011000000000 : n22046_o;
  assign n22059_o = n20500_o[3:2];
  /* loadstore1.vhdl:859:13  */
  assign n22060_o = n22011_o ? n22059_o : n22048_o;
  assign n22061_o = n20500_o[12];
  /* loadstore1.vhdl:859:13  */
  assign n22062_o = n22011_o ? n22061_o : n22050_o;
  assign n22063_o = n20500_o[14];
  /* loadstore1.vhdl:859:13  */
  assign n22064_o = n22011_o ? n22063_o : n22052_o;
  assign n22065_o = {n22057_o, n22054_o};
  assign n22066_o = {n22009_o, n22058_o};
  /* loadstore1.vhdl:857:9  */
  assign n22067_o = n21966_o ? n22065_o : n21934_o;
  /* loadstore1.vhdl:857:9  */
  assign n22068_o = n21966_o ? n22066_o : n22007_o;
  assign n22069_o = n20500_o[3:2];
  /* loadstore1.vhdl:857:9  */
  assign n22070_o = n21966_o ? n22060_o : n22069_o;
  assign n22071_o = n20500_o[12];
  /* loadstore1.vhdl:857:9  */
  assign n22072_o = n21966_o ? n22062_o : n22071_o;
  assign n22073_o = n20500_o[14];
  /* loadstore1.vhdl:857:9  */
  assign n22074_o = n21966_o ? n22064_o : n22073_o;
  assign n22076_o = n20500_o[1:0];
  assign n22078_o = n20500_o[11:4];
  assign n22079_o = n20500_o[15];
  assign n22080_o = n20500_o[13];
  /* loadstore1.vhdl:883:17  */
  assign n22081_o = r2[309:308];
  /* loadstore1.vhdl:884:9  */
  assign n22083_o = n22081_o == 2'b00;
  /* loadstore1.vhdl:889:30  */
  assign n22084_o = r2[373:310];
  /* loadstore1.vhdl:887:9  */
  assign n22086_o = n22081_o == 2'b01;
  /* loadstore1.vhdl:890:9  */
  assign n22088_o = n22081_o == 2'b10;
  assign n22089_o = {n21047_o, n21009_o, n20971_o, n20933_o, n20895_o, n20857_o, n20819_o, n20781_o};
  assign n22090_o = {n22088_o, n22086_o, n22083_o};
  /* loadstore1.vhdl:883:9  */
  always @*
    case (n22090_o)
      3'b100: n22091_o = load_dp_data;
      3'b010: n22091_o = n22084_o;
      3'b001: n22091_o = n21759_o;
      default: n22091_o = n22089_o;
    endcase
  /* loadstore1.vhdl:901:38  */
  assign n22092_o = stage1_req[2];
  /* loadstore1.vhdl:902:38  */
  assign n22093_o = stage1_req[5];
  /* loadstore1.vhdl:903:36  */
  assign n22094_o = stage1_req[191];
  /* loadstore1.vhdl:904:41  */
  assign n22095_o = stage1_req[187];
  /* loadstore1.vhdl:905:40  */
  assign n22096_o = stage1_req[188];
  /* loadstore1.vhdl:906:45  */
  assign n22097_o = stage1_req[189];
  /* loadstore1.vhdl:907:38  */
  assign n22098_o = stage1_req[77:14];
  /* loadstore1.vhdl:908:42  */
  assign n22099_o = stage1_req[85:78];
  /* loadstore1.vhdl:909:43  */
  assign n22100_o = stage1_req[192];
  /* loadstore1.vhdl:910:43  */
  assign n22101_o = stage1_req[193];
  /* loadstore1.vhdl:913:30  */
  assign n22102_o = r2[272:0];
  /* loadstore1.vhdl:913:34  */
  assign n22103_o = n22102_o[2];
  /* loadstore1.vhdl:914:30  */
  assign n22104_o = r2[272:0];
  /* loadstore1.vhdl:914:34  */
  assign n22105_o = n22104_o[5];
  /* loadstore1.vhdl:915:28  */
  assign n22106_o = r2[272:0];
  /* loadstore1.vhdl:915:32  */
  assign n22107_o = n22106_o[191];
  /* loadstore1.vhdl:916:33  */
  assign n22108_o = r2[272:0];
  /* loadstore1.vhdl:916:37  */
  assign n22109_o = n22108_o[187];
  /* loadstore1.vhdl:917:32  */
  assign n22110_o = r2[272:0];
  /* loadstore1.vhdl:917:36  */
  assign n22111_o = n22110_o[188];
  /* loadstore1.vhdl:918:37  */
  assign n22112_o = r2[272:0];
  /* loadstore1.vhdl:918:41  */
  assign n22113_o = n22112_o[189];
  /* loadstore1.vhdl:919:30  */
  assign n22114_o = r2[272:0];
  /* loadstore1.vhdl:919:34  */
  assign n22115_o = n22114_o[77:14];
  /* loadstore1.vhdl:920:34  */
  assign n22116_o = r2[272:0];
  /* loadstore1.vhdl:920:38  */
  assign n22117_o = n22116_o[85:78];
  /* loadstore1.vhdl:921:35  */
  assign n22118_o = r2[272:0];
  /* loadstore1.vhdl:921:39  */
  assign n22119_o = n22118_o[192];
  /* loadstore1.vhdl:922:35  */
  assign n22120_o = r2[272:0];
  /* loadstore1.vhdl:922:39  */
  assign n22121_o = n22120_o[193];
  assign n22122_o = {n22115_o, n22121_o, n22119_o, n22113_o, n22111_o, n22109_o, n22107_o, n22105_o, n22103_o};
  assign n22123_o = {n22098_o, n22101_o, n22100_o, n22097_o, n22096_o, n22095_o, n22094_o, n22093_o, n22092_o};
  /* loadstore1.vhdl:899:9  */
  assign n22124_o = stage1_issue_enable ? stage1_dcreq : n21946_o;
  /* loadstore1.vhdl:899:9  */
  assign n22125_o = stage1_issue_enable ? n22123_o : n22122_o;
  /* loadstore1.vhdl:899:9  */
  assign n22126_o = stage1_issue_enable ? n22099_o : n22117_o;
  /* loadstore1.vhdl:927:30  */
  assign n22127_o = r2[272:0];
  /* loadstore1.vhdl:927:34  */
  assign n22128_o = n22127_o[157:94];
  /* loadstore1.vhdl:924:9  */
  assign n22129_o = stage1_dreq ? store_data : n22128_o;
  /* loadstore1.vhdl:929:26  */
  assign n22130_o = r2[272:0];
  /* loadstore1.vhdl:929:30  */
  assign n22131_o = n22130_o[0];
  /* loadstore1.vhdl:929:43  */
  assign n22132_o = r2[272:0];
  /* loadstore1.vhdl:929:47  */
  assign n22133_o = n22132_o[194];
  /* loadstore1.vhdl:929:36  */
  assign n22134_o = n22131_o & n22133_o;
  /* loadstore1.vhdl:929:64  */
  assign n22135_o = n19358_o[0];
  /* loadstore1.vhdl:929:55  */
  assign n22136_o = n22134_o & n22135_o;
  /* loadstore1.vhdl:933:27  */
  assign n22137_o = r2[272:0];
  /* loadstore1.vhdl:933:31  */
  assign n22138_o = n22137_o[9];
  /* loadstore1.vhdl:934:26  */
  assign n22139_o = r2[272:0];
  /* loadstore1.vhdl:934:30  */
  assign n22140_o = n22139_o[2];
  /* loadstore1.vhdl:935:26  */
  assign n22141_o = r2[272:0];
  /* loadstore1.vhdl:935:30  */
  assign n22142_o = n22141_o[193];
  /* loadstore1.vhdl:936:27  */
  assign n22143_o = r2[272:0];
  /* loadstore1.vhdl:936:31  */
  assign n22144_o = n22143_o[4];
  /* loadstore1.vhdl:938:26  */
  assign n22145_o = r2[272:0];
  /* loadstore1.vhdl:938:30  */
  assign n22146_o = n22145_o[204:195];
  /* loadstore1.vhdl:939:26  */
  assign n22147_o = r2[272:0];
  /* loadstore1.vhdl:939:30  */
  assign n22148_o = n22147_o[77:14];
  /* loadstore1.vhdl:940:27  */
  assign n22149_o = r2[272:0];
  /* loadstore1.vhdl:940:31  */
  assign n22150_o = n22149_o[205];
  /* loadstore1.vhdl:941:24  */
  assign n22151_o = r2[272:0];
  /* loadstore1.vhdl:941:28  */
  assign n22152_o = n22151_o[157:94];
  /* loadstore1.vhdl:945:31  */
  assign n22153_o = r2[272:0];
  /* loadstore1.vhdl:945:35  */
  assign n22154_o = n22153_o[160:158];
  /* loadstore1.vhdl:946:44  */
  assign n22155_o = n21958_o | n21960_o;
  /* loadstore1.vhdl:947:31  */
  assign n22156_o = r2[272:0];
  /* loadstore1.vhdl:947:35  */
  assign n22157_o = n22156_o[167:161];
  /* loadstore1.vhdl:949:26  */
  assign n22158_o = r2[272:0];
  /* loadstore1.vhdl:949:30  */
  assign n22159_o = n22158_o[186:182];
  /* loadstore1.vhdl:950:24  */
  assign n22160_o = r2[272:0];
  /* loadstore1.vhdl:950:28  */
  assign n22161_o = n22160_o[190];
  /* loadstore1.vhdl:950:31  */
  assign n22162_o = n22161_o & complete;
  /* loadstore1.vhdl:951:34  */
  assign n22163_o = n19358_o[65];
  /* loadstore1.vhdl:952:31  */
  assign n22164_o = r3[285];
  /* loadstore1.vhdl:953:30  */
  assign n22165_o = r3[297:286];
  /* loadstore1.vhdl:954:26  */
  assign n22166_o = r3[361:298];
  /* loadstore1.vhdl:955:26  */
  assign n22167_o = r3[377:362];
  /* loadstore1.vhdl:960:31  */
  assign n22168_o = r3[285];
  /* loadstore1.vhdl:962:22  */
  assign n22169_o = r3[380:378];
  /* loadstore1.vhdl:965:32  */
  assign n22170_o = r2[272:0];
  /* loadstore1.vhdl:965:36  */
  assign n22171_o = n22170_o[0];
  /* loadstore1.vhdl:965:60  */
  assign n22172_o = complete | n21963_o;
  /* loadstore1.vhdl:965:73  */
  assign n22173_o = n22172_o | n21966_o;
  /* loadstore1.vhdl:965:46  */
  assign n22174_o = ~n22173_o;
  /* loadstore1.vhdl:965:42  */
  assign n22175_o = n22171_o & n22174_o;
  assign n22176_o = {n21940_o, n22006_o, n21999_o, n22079_o, n22074_o, n22080_o, n22072_o, n22078_o, n22070_o, n22076_o, n22068_o, n21966_o, n21996_o, n21701_o, n21054_o, n21049_o, n22067_o, n21710_o, n21932_o, n21941_o, n21995_o};
  /* loadstore1.vhdl:275:9  */
  always @(posedge clk)
    n22184_q <= n19449_o;
  /* loadstore1.vhdl:275:9  */
  always @(posedge clk)
    n22185_q <= n19451_o;
  /* loadstore1.vhdl:275:9  */
  always @(posedge clk)
    n22186_q <= n19453_o;
  /* loadstore1.vhdl:275:9  */
  always @(posedge clk)
    n22187_q <= n19443_o;
  /* loadstore1.vhdl:275:9  */
  assign n22188_o = {n19462_o, n19541_o, n19538_o};
  assign n22189_o = {n19585_o, n19581_o, n19639_o, 29'b00000000000000000000000000000};
  assign n22190_o = {n22308_o, n22294_o, n22280_o, n22266_o, n22252_o, n22238_o, n22224_o, n22210_o};
  /* loadstore1.vhdl:275:9  */
  always @(posedge clk)
    n22191_q <= stage1_dcreq;
  /* loadstore1.vhdl:275:9  */
  assign n22192_o = {n22168_o, in_progress, busy};
  assign n22193_o = {n22167_o, n22166_o, n22165_o, n22164_o, n22163_o, n22162_o, n22159_o, n22091_o, n22157_o, n22155_o, n22154_o, complete};
  assign n22194_o = {n22126_o, n22129_o, n22125_o, n22136_o, n22124_o};
  assign n22195_o = {n22152_o, n22148_o, n22146_o, n22142_o, n22140_o, n22138_o, n21954_o, n22150_o, n22144_o, n21950_o};
  assign n22197_o = r1[101:94];
  /* loadstore1.vhdl:38:9  */
  assign n22198_o = r1[109:102];
  /* loadstore1.vhdl:36:9  */
  assign n22199_o = r1[117:110];
  /* loadstore1.vhdl:31:9  */
  assign n22200_o = r1[125:118];
  /* loadstore1.vhdl:28:9  */
  assign n22201_o = r1[133:126];
  /* loadstore1.vhdl:26:9  */
  assign n22202_o = r1[141:134];
  /* loadstore1.vhdl:25:9  */
  assign n22203_o = r1[149:142];
  assign n22204_o = r1[157:150];
  /* loadstore1.vhdl:595:68  */
  assign n22205_o = n20182_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22205_o)
      2'b00: n22206_o = n22197_o;
      2'b01: n22206_o = n22198_o;
      2'b10: n22206_o = n22199_o;
      2'b11: n22206_o = n22200_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22207_o = n20182_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22207_o)
      2'b00: n22208_o = n22201_o;
      2'b01: n22208_o = n22202_o;
      2'b10: n22208_o = n22203_o;
      2'b11: n22208_o = n22204_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22209_o = n20182_o[2];
  /* loadstore1.vhdl:595:68  */
  assign n22210_o = n22209_o ? n22208_o : n22206_o;
  /* loadstore1.vhdl:595:68  */
  assign n22211_o = r1[101:94];
  /* loadstore1.vhdl:595:68  */
  assign n22212_o = r1[109:102];
  assign n22213_o = r1[117:110];
  assign n22214_o = r1[125:118];
  assign n22215_o = r1[133:126];
  assign n22216_o = r1[141:134];
  assign n22217_o = r1[149:142];
  assign n22218_o = r1[157:150];
  /* loadstore1.vhdl:595:68  */
  assign n22219_o = n20195_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22219_o)
      2'b00: n22220_o = n22211_o;
      2'b01: n22220_o = n22212_o;
      2'b10: n22220_o = n22213_o;
      2'b11: n22220_o = n22214_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22221_o = n20195_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22221_o)
      2'b00: n22222_o = n22215_o;
      2'b01: n22222_o = n22216_o;
      2'b10: n22222_o = n22217_o;
      2'b11: n22222_o = n22218_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22223_o = n20195_o[2];
  /* loadstore1.vhdl:595:68  */
  assign n22224_o = n22223_o ? n22222_o : n22220_o;
  /* loadstore1.vhdl:595:68  */
  assign n22225_o = r1[101:94];
  /* loadstore1.vhdl:595:68  */
  assign n22226_o = r1[109:102];
  assign n22227_o = r1[117:110];
  assign n22228_o = r1[125:118];
  assign n22229_o = r1[133:126];
  assign n22230_o = r1[141:134];
  assign n22231_o = r1[149:142];
  assign n22232_o = r1[157:150];
  /* loadstore1.vhdl:595:68  */
  assign n22233_o = n20208_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22233_o)
      2'b00: n22234_o = n22225_o;
      2'b01: n22234_o = n22226_o;
      2'b10: n22234_o = n22227_o;
      2'b11: n22234_o = n22228_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22235_o = n20208_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22235_o)
      2'b00: n22236_o = n22229_o;
      2'b01: n22236_o = n22230_o;
      2'b10: n22236_o = n22231_o;
      2'b11: n22236_o = n22232_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22237_o = n20208_o[2];
  /* loadstore1.vhdl:595:68  */
  assign n22238_o = n22237_o ? n22236_o : n22234_o;
  /* loadstore1.vhdl:595:68  */
  assign n22239_o = r1[101:94];
  /* loadstore1.vhdl:595:68  */
  assign n22240_o = r1[109:102];
  assign n22241_o = r1[117:110];
  assign n22242_o = r1[125:118];
  assign n22243_o = r1[133:126];
  assign n22244_o = r1[141:134];
  assign n22245_o = r1[149:142];
  assign n22246_o = r1[157:150];
  /* loadstore1.vhdl:595:68  */
  assign n22247_o = n20221_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22247_o)
      2'b00: n22248_o = n22239_o;
      2'b01: n22248_o = n22240_o;
      2'b10: n22248_o = n22241_o;
      2'b11: n22248_o = n22242_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22249_o = n20221_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22249_o)
      2'b00: n22250_o = n22243_o;
      2'b01: n22250_o = n22244_o;
      2'b10: n22250_o = n22245_o;
      2'b11: n22250_o = n22246_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22251_o = n20221_o[2];
  /* loadstore1.vhdl:595:68  */
  assign n22252_o = n22251_o ? n22250_o : n22248_o;
  /* loadstore1.vhdl:595:68  */
  assign n22253_o = r1[101:94];
  /* loadstore1.vhdl:595:68  */
  assign n22254_o = r1[109:102];
  assign n22255_o = r1[117:110];
  assign n22256_o = r1[125:118];
  /* helpers.vhdl:237:18  */
  assign n22257_o = r1[133:126];
  assign n22258_o = r1[141:134];
  /* helpers.vhdl:236:18  */
  assign n22259_o = r1[149:142];
  assign n22260_o = r1[157:150];
  /* loadstore1.vhdl:595:68  */
  assign n22261_o = n20234_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22261_o)
      2'b00: n22262_o = n22253_o;
      2'b01: n22262_o = n22254_o;
      2'b10: n22262_o = n22255_o;
      2'b11: n22262_o = n22256_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22263_o = n20234_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22263_o)
      2'b00: n22264_o = n22257_o;
      2'b01: n22264_o = n22258_o;
      2'b10: n22264_o = n22259_o;
      2'b11: n22264_o = n22260_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22265_o = n20234_o[2];
  /* loadstore1.vhdl:595:68  */
  assign n22266_o = n22265_o ? n22264_o : n22262_o;
  /* loadstore1.vhdl:595:68  */
  assign n22267_o = r1[101:94];
  /* loadstore1.vhdl:595:68  */
  assign n22268_o = r1[109:102];
  assign n22269_o = r1[117:110];
  /* helpers.vhdl:30:14  */
  assign n22270_o = r1[125:118];
  assign n22271_o = r1[133:126];
  assign n22272_o = r1[141:134];
  assign n22273_o = r1[149:142];
  assign n22274_o = r1[157:150];
  /* loadstore1.vhdl:595:68  */
  assign n22275_o = n20247_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22275_o)
      2'b00: n22276_o = n22267_o;
      2'b01: n22276_o = n22268_o;
      2'b10: n22276_o = n22269_o;
      2'b11: n22276_o = n22270_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22277_o = n20247_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22277_o)
      2'b00: n22278_o = n22271_o;
      2'b01: n22278_o = n22272_o;
      2'b10: n22278_o = n22273_o;
      2'b11: n22278_o = n22274_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22279_o = n20247_o[2];
  /* loadstore1.vhdl:595:68  */
  assign n22280_o = n22279_o ? n22278_o : n22276_o;
  /* loadstore1.vhdl:595:68  */
  assign n22281_o = r1[101:94];
  /* loadstore1.vhdl:595:68  */
  assign n22282_o = r1[109:102];
  assign n22283_o = r1[117:110];
  assign n22284_o = r1[125:118];
  assign n22285_o = r1[133:126];
  /* helpers.vhdl:259:18  */
  assign n22286_o = r1[141:134];
  assign n22287_o = r1[149:142];
  /* helpers.vhdl:258:18  */
  assign n22288_o = r1[157:150];
  /* loadstore1.vhdl:595:68  */
  assign n22289_o = n20260_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22289_o)
      2'b00: n22290_o = n22281_o;
      2'b01: n22290_o = n22282_o;
      2'b10: n22290_o = n22283_o;
      2'b11: n22290_o = n22284_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22291_o = n20260_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22291_o)
      2'b00: n22292_o = n22285_o;
      2'b01: n22292_o = n22286_o;
      2'b10: n22292_o = n22287_o;
      2'b11: n22292_o = n22288_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22293_o = n20260_o[2];
  /* loadstore1.vhdl:595:68  */
  assign n22294_o = n22293_o ? n22292_o : n22290_o;
  /* loadstore1.vhdl:595:68  */
  assign n22295_o = r1[101:94];
  /* loadstore1.vhdl:595:68  */
  assign n22296_o = r1[109:102];
  /* helpers.vhdl:31:14  */
  assign n22297_o = r1[117:110];
  assign n22298_o = r1[125:118];
  /* helpers.vhdl:31:14  */
  assign n22299_o = r1[133:126];
  assign n22300_o = r1[141:134];
  assign n22301_o = r1[149:142];
  assign n22302_o = r1[157:150];
  /* loadstore1.vhdl:595:68  */
  assign n22303_o = n20273_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22303_o)
      2'b00: n22304_o = n22295_o;
      2'b01: n22304_o = n22296_o;
      2'b10: n22304_o = n22297_o;
      2'b11: n22304_o = n22298_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22305_o = n20273_o[1:0];
  /* loadstore1.vhdl:595:68  */
  always @*
    case (n22305_o)
      2'b00: n22306_o = n22299_o;
      2'b01: n22306_o = n22300_o;
      2'b10: n22306_o = n22301_o;
      2'b11: n22306_o = n22302_o;
    endcase
  /* loadstore1.vhdl:595:68  */
  assign n22307_o = n20273_o[2];
  /* loadstore1.vhdl:595:68  */
  assign n22308_o = n22307_o ? n22306_o : n22304_o;
  /* loadstore1.vhdl:595:68  */
  assign n22309_o = n19358_o[8:1];
  /* loadstore1.vhdl:595:68  */
  assign n22310_o = n19358_o[16:9];
  /* helpers.vhdl:279:18  */
  assign n22311_o = n19358_o[24:17];
  assign n22312_o = n19358_o[32:25];
  /* helpers.vhdl:278:18  */
  assign n22313_o = n19358_o[40:33];
  assign n22314_o = n19358_o[48:41];
  /* helpers.vhdl:277:18  */
  assign n22315_o = n19358_o[56:49];
  assign n22316_o = n19358_o[64:57];
  /* loadstore1.vhdl:685:63  */
  assign n22317_o = n20504_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22317_o)
      2'b00: n22318_o = n22309_o;
      2'b01: n22318_o = n22310_o;
      2'b10: n22318_o = n22311_o;
      2'b11: n22318_o = n22312_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22319_o = n20504_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22319_o)
      2'b00: n22320_o = n22313_o;
      2'b01: n22320_o = n22314_o;
      2'b10: n22320_o = n22315_o;
      2'b11: n22320_o = n22316_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22321_o = n20504_o[2];
  /* loadstore1.vhdl:685:63  */
  assign n22322_o = n22321_o ? n22320_o : n22318_o;
  /* loadstore1.vhdl:685:63  */
  assign n22323_o = n19358_o[8:1];
  /* loadstore1.vhdl:685:63  */
  assign n22324_o = n19358_o[16:9];
  assign n22325_o = n19358_o[24:17];
  assign n22326_o = n19358_o[32:25];
  assign n22327_o = n19358_o[40:33];
  assign n22328_o = n19358_o[48:41];
  assign n22329_o = n19358_o[56:49];
  assign n22330_o = n19358_o[64:57];
  /* loadstore1.vhdl:685:63  */
  assign n22331_o = n20513_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22331_o)
      2'b00: n22332_o = n22323_o;
      2'b01: n22332_o = n22324_o;
      2'b10: n22332_o = n22325_o;
      2'b11: n22332_o = n22326_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22333_o = n20513_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22333_o)
      2'b00: n22334_o = n22327_o;
      2'b01: n22334_o = n22328_o;
      2'b10: n22334_o = n22329_o;
      2'b11: n22334_o = n22330_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22335_o = n20513_o[2];
  /* loadstore1.vhdl:685:63  */
  assign n22336_o = n22335_o ? n22334_o : n22332_o;
  /* loadstore1.vhdl:685:63  */
  assign n22337_o = n19358_o[8:1];
  /* loadstore1.vhdl:685:63  */
  assign n22338_o = n19358_o[16:9];
  assign n22339_o = n19358_o[24:17];
  assign n22340_o = n19358_o[32:25];
  assign n22341_o = n19358_o[40:33];
  assign n22342_o = n19358_o[48:41];
  assign n22343_o = n19358_o[56:49];
  assign n22344_o = n19358_o[64:57];
  /* loadstore1.vhdl:685:63  */
  assign n22345_o = n20522_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22345_o)
      2'b00: n22346_o = n22337_o;
      2'b01: n22346_o = n22338_o;
      2'b10: n22346_o = n22339_o;
      2'b11: n22346_o = n22340_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22347_o = n20522_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22347_o)
      2'b00: n22348_o = n22341_o;
      2'b01: n22348_o = n22342_o;
      2'b10: n22348_o = n22343_o;
      2'b11: n22348_o = n22344_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22349_o = n20522_o[2];
  /* loadstore1.vhdl:685:63  */
  assign n22350_o = n22349_o ? n22348_o : n22346_o;
  /* loadstore1.vhdl:685:63  */
  assign n22351_o = n19358_o[8:1];
  /* loadstore1.vhdl:685:63  */
  assign n22352_o = n19358_o[16:9];
  /* helpers.vhdl:29:14  */
  assign n22353_o = n19358_o[24:17];
  /* helpers.vhdl:29:14  */
  assign n22354_o = n19358_o[32:25];
  assign n22355_o = n19358_o[40:33];
  /* helpers.vhdl:29:14  */
  assign n22356_o = n19358_o[48:41];
  /* helpers.vhdl:292:18  */
  assign n22357_o = n19358_o[56:49];
  assign n22358_o = n19358_o[64:57];
  /* loadstore1.vhdl:685:63  */
  assign n22359_o = n20531_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22359_o)
      2'b00: n22360_o = n22351_o;
      2'b01: n22360_o = n22352_o;
      2'b10: n22360_o = n22353_o;
      2'b11: n22360_o = n22354_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22361_o = n20531_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22361_o)
      2'b00: n22362_o = n22355_o;
      2'b01: n22362_o = n22356_o;
      2'b10: n22362_o = n22357_o;
      2'b11: n22362_o = n22358_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22363_o = n20531_o[2];
  /* loadstore1.vhdl:685:63  */
  assign n22364_o = n22363_o ? n22362_o : n22360_o;
  /* loadstore1.vhdl:685:63  */
  assign n22365_o = n19358_o[8:1];
  /* loadstore1.vhdl:685:63  */
  assign n22366_o = n19358_o[16:9];
  assign n22367_o = n19358_o[24:17];
  /* loadstore1.vhdl:685:66  */
  assign n22368_o = n19358_o[32:25];
  assign n22369_o = n19358_o[40:33];
  /* loadstore1.vhdl:684:47  */
  assign n22370_o = n19358_o[48:41];
  assign n22371_o = n19358_o[56:49];
  /* loadstore1.vhdl:684:47  */
  assign n22372_o = n19358_o[64:57];
  /* loadstore1.vhdl:685:63  */
  assign n22373_o = n20540_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22373_o)
      2'b00: n22374_o = n22365_o;
      2'b01: n22374_o = n22366_o;
      2'b10: n22374_o = n22367_o;
      2'b11: n22374_o = n22368_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22375_o = n20540_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22375_o)
      2'b00: n22376_o = n22369_o;
      2'b01: n22376_o = n22370_o;
      2'b10: n22376_o = n22371_o;
      2'b11: n22376_o = n22372_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22377_o = n20540_o[2];
  /* loadstore1.vhdl:685:63  */
  assign n22378_o = n22377_o ? n22376_o : n22374_o;
  /* loadstore1.vhdl:685:63  */
  assign n22379_o = n19358_o[8:1];
  /* loadstore1.vhdl:685:63  */
  assign n22380_o = n19358_o[16:9];
  /* loadstore1.vhdl:684:18  */
  assign n22381_o = n19358_o[24:17];
  /* loadstore1.vhdl:685:66  */
  assign n22382_o = n19358_o[32:25];
  assign n22383_o = n19358_o[40:33];
  /* loadstore1.vhdl:684:47  */
  assign n22384_o = n19358_o[48:41];
  assign n22385_o = n19358_o[56:49];
  /* loadstore1.vhdl:684:47  */
  assign n22386_o = n19358_o[64:57];
  /* loadstore1.vhdl:685:63  */
  assign n22387_o = n20549_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22387_o)
      2'b00: n22388_o = n22379_o;
      2'b01: n22388_o = n22380_o;
      2'b10: n22388_o = n22381_o;
      2'b11: n22388_o = n22382_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22389_o = n20549_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22389_o)
      2'b00: n22390_o = n22383_o;
      2'b01: n22390_o = n22384_o;
      2'b10: n22390_o = n22385_o;
      2'b11: n22390_o = n22386_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22391_o = n20549_o[2];
  /* loadstore1.vhdl:685:63  */
  assign n22392_o = n22391_o ? n22390_o : n22388_o;
  /* loadstore1.vhdl:685:63  */
  assign n22393_o = n19358_o[8:1];
  /* loadstore1.vhdl:685:63  */
  assign n22394_o = n19358_o[16:9];
  /* loadstore1.vhdl:684:18  */
  assign n22395_o = n19358_o[24:17];
  /* loadstore1.vhdl:685:66  */
  assign n22396_o = n19358_o[32:25];
  assign n22397_o = n19358_o[40:33];
  /* loadstore1.vhdl:684:47  */
  assign n22398_o = n19358_o[48:41];
  assign n22399_o = n19358_o[56:49];
  /* loadstore1.vhdl:684:47  */
  assign n22400_o = n19358_o[64:57];
  /* loadstore1.vhdl:685:63  */
  assign n22401_o = n20558_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22401_o)
      2'b00: n22402_o = n22393_o;
      2'b01: n22402_o = n22394_o;
      2'b10: n22402_o = n22395_o;
      2'b11: n22402_o = n22396_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22403_o = n20558_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22403_o)
      2'b00: n22404_o = n22397_o;
      2'b01: n22404_o = n22398_o;
      2'b10: n22404_o = n22399_o;
      2'b11: n22404_o = n22400_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22405_o = n20558_o[2];
  /* loadstore1.vhdl:685:63  */
  assign n22406_o = n22405_o ? n22404_o : n22402_o;
  /* loadstore1.vhdl:685:63  */
  assign n22407_o = n19358_o[8:1];
  /* loadstore1.vhdl:685:63  */
  assign n22408_o = n19358_o[16:9];
  /* loadstore1.vhdl:684:18  */
  assign n22409_o = n19358_o[24:17];
  /* loadstore1.vhdl:685:66  */
  assign n22410_o = n19358_o[32:25];
  assign n22411_o = n19358_o[40:33];
  /* loadstore1.vhdl:684:47  */
  assign n22412_o = n19358_o[48:41];
  assign n22413_o = n19358_o[56:49];
  /* loadstore1.vhdl:684:47  */
  assign n22414_o = n19358_o[64:57];
  /* loadstore1.vhdl:685:63  */
  assign n22415_o = n20567_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22415_o)
      2'b00: n22416_o = n22407_o;
      2'b01: n22416_o = n22408_o;
      2'b10: n22416_o = n22409_o;
      2'b11: n22416_o = n22410_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22417_o = n20567_o[1:0];
  /* loadstore1.vhdl:685:63  */
  always @*
    case (n22417_o)
      2'b00: n22418_o = n22411_o;
      2'b01: n22418_o = n22412_o;
      2'b10: n22418_o = n22413_o;
      2'b11: n22418_o = n22414_o;
    endcase
  /* loadstore1.vhdl:685:63  */
  assign n22419_o = n20567_o[2];
  /* loadstore1.vhdl:685:63  */
  assign n22420_o = n22419_o ? n22418_o : n22416_o;
endmodule

module fpu
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  clk,
   input  rst,
   input  e_in_valid,
   input  [5:0] e_in_op,
   input  [63:0] e_in_nia,
   input  [2:0] e_in_itag,
   input  [31:0] e_in_insn,
   input  e_in_single,
   input  [1:0] e_in_fe_mode,
   input  [63:0] e_in_fra,
   input  [63:0] e_in_frb,
   input  [63:0] e_in_frc,
   input  [6:0] e_in_frt,
   input  e_in_rc,
   input  e_in_out_cr,
   output e_out_busy,
   output e_out_exception,
   output w_out_valid,
   output w_out_interrupt,
   output [2:0] w_out_instr_tag,
   output w_out_write_enable,
   output [6:0] w_out_write_reg,
   output [63:0] w_out_write_data,
   output w_out_write_cr_enable,
   output [7:0] w_out_write_cr_mask,
   output [31:0] w_out_write_cr_data,
   output [11:0] w_out_intr_vec,
   output [63:0] w_out_srr0,
   output [15:0] w_out_srr1);
  wire [309:0] n12968_o;
  wire n12970_o;
  wire n12971_o;
  wire n12973_o;
  wire n12974_o;
  wire [2:0] n12975_o;
  wire n12976_o;
  wire [6:0] n12977_o;
  wire [63:0] n12978_o;
  wire n12979_o;
  wire [7:0] n12980_o;
  wire [31:0] n12981_o;
  wire [11:0] n12982_o;
  wire [63:0] n12983_o;
  wire [15:0] n12984_o;
  wire [721:0] r;
  wire [721:0] rin;
  wire [63:0] fp_result;
  wire [1:0] opsel_b;
  wire [1:0] opsel_r;
  wire [1:0] opsel_s;
  wire opsel_ainv;
  wire opsel_mask;
  wire opsel_binv;
  wire [63:0] in_a;
  wire [63:0] in_b;
  wire [63:0] result;
  wire carry_in;
  wire r_hi_nz;
  wire r_lo_nz;
  wire s_nz;
  wire [3:0] misc_sel;
  wire [258:0] f_to_multiply;
  wire [129:0] multiply_to_f;
  wire [1:0] msel_1;
  wire [1:0] msel_2;
  wire [1:0] msel_add;
  wire msel_inv;
  wire [18:0] inverse_est;
  wire fpu_multiply_0_m_out_valid;
  wire [127:0] fpu_multiply_0_m_out_result;
  wire fpu_multiply_0_m_out_overflow;
  wire n12985_o;
  wire [63:0] n12986_o;
  wire [63:0] n12987_o;
  wire [127:0] n12988_o;
  wire n12989_o;
  wire n12990_o;
  wire [129:0] n12991_o;
  wire [9:0] n13001_o;
  wire [9:0] n13002_o;
  wire [9:0] n13003_o;
  wire [116:0] n13004_o;
  wire [116:0] n13005_o;
  wire [116:0] n13006_o;
  wire [31:0] n13007_o;
  wire [31:0] n13008_o;
  wire [517:0] n13009_o;
  wire [517:0] n13010_o;
  wire [517:0] n13011_o;
  wire n13012_o;
  wire n13013_o;
  wire [43:0] n13014_o;
  wire [43:0] n13015_o;
  wire [43:0] n13016_o;
  wire [721:0] n13017_o;
  wire n13024_o;
  wire [1:0] n13025_o;
  wire [1:0] n13027_o;
  wire [7:0] n13028_o;
  wire [9:0] n13029_o;
  wire [9:0] n13032_o;
  wire [18:0] n13037_o;
  wire n13042_o;
  wire n13043_o;
  wire n13044_o;
  wire n13045_o;
  wire n13046_o;
  wire n13047_o;
  wire [2:0] n13048_o;
  wire n13049_o;
  wire [6:0] n13050_o;
  wire n13051_o;
  wire n13052_o;
  wire n13053_o;
  wire n13054_o;
  wire n13055_o;
  wire [7:0] n13056_o;
  wire [3:0] n13057_o;
  wire [3:0] n13058_o;
  wire [7:0] n13059_o;
  wire [3:0] n13060_o;
  wire [11:0] n13061_o;
  wire [3:0] n13062_o;
  wire [15:0] n13063_o;
  wire [3:0] n13064_o;
  wire [19:0] n13065_o;
  wire [3:0] n13066_o;
  wire [23:0] n13067_o;
  wire [3:0] n13068_o;
  wire [27:0] n13069_o;
  wire [3:0] n13070_o;
  wire [31:0] n13071_o;
  wire n13072_o;
  wire [63:0] n13074_o;
  wire n13075_o;
  wire n13076_o;
  wire n13077_o;
  wire [3:0] n13092_o;
  wire [3:0] n13093_o;
  wire [3:0] n13094_o;
  wire [3:0] n13095_o;
  wire [15:0] n13096_o;
  wire [6:0] n13151_o;
  wire n13152_o;
  wire [31:0] n13153_o;
  wire [63:0] n13154_o;
  wire [5:0] n13155_o;
  wire [2:0] n13156_o;
  wire [1:0] n13157_o;
  wire n13158_o;
  wire [6:0] n13159_o;
  wire n13160_o;
  wire n13161_o;
  wire n13163_o;
  wire n13164_o;
  wire n13165_o;
  wire n13166_o;
  wire [31:0] n13171_o;
  wire [2:0] n13176_o;
  wire n13184_o;
  wire n13187_o;
  wire n13190_o;
  wire n13193_o;
  wire n13196_o;
  wire n13199_o;
  wire n13202_o;
  wire n13205_o;
  wire [7:0] n13207_o;
  reg [7:0] n13208_o;
  wire [7:0] n13209_o;
  wire [5:0] n13210_o;
  wire n13212_o;
  wire n13215_o;
  wire [1:0] n13220_o;
  wire [2:0] n13222_o;
  wire [63:0] n13229_o;
  wire n13239_o;
  wire [10:0] n13243_o;
  wire n13244_o;
  wire [10:0] n13246_o;
  wire n13247_o;
  wire [51:0] n13249_o;
  wire n13250_o;
  wire n13252_o;
  wire [10:0] n13253_o;
  wire [12:0] n13254_o;
  wire [12:0] n13256_o;
  wire n13257_o;
  wire [12:0] n13259_o;
  wire [9:0] n13261_o;
  wire [51:0] n13262_o;
  wire [61:0] n13263_o;
  wire [63:0] n13265_o;
  wire [1:0] n13266_o;
  wire [2:0] n13267_o;
  wire n13270_o;
  wire n13273_o;
  wire n13276_o;
  wire n13279_o;
  wire n13282_o;
  wire [4:0] n13284_o;
  reg [1:0] n13285_o;
  wire n13287_o;
  wire n13288_o;
  wire n13289_o;
  wire [1:0] n13292_o;
  wire [76:0] n13293_o;
  wire [76:0] n13294_o;
  wire [1:0] n13295_o;
  wire [76:0] n13296_o;
  wire [79:0] n13300_o;
  wire [63:0] n13302_o;
  wire n13312_o;
  wire [10:0] n13316_o;
  wire n13317_o;
  wire [10:0] n13319_o;
  wire n13320_o;
  wire [51:0] n13322_o;
  wire n13323_o;
  wire n13325_o;
  wire [10:0] n13326_o;
  wire [12:0] n13327_o;
  wire [12:0] n13329_o;
  wire n13330_o;
  wire [12:0] n13332_o;
  wire [9:0] n13334_o;
  wire [51:0] n13335_o;
  wire [61:0] n13336_o;
  wire [63:0] n13338_o;
  wire [1:0] n13339_o;
  wire [2:0] n13340_o;
  wire n13343_o;
  wire n13346_o;
  wire n13349_o;
  wire n13352_o;
  wire n13355_o;
  wire [4:0] n13357_o;
  reg [1:0] n13358_o;
  wire n13360_o;
  wire n13361_o;
  wire n13362_o;
  wire [1:0] n13365_o;
  wire [76:0] n13366_o;
  wire [76:0] n13367_o;
  wire [1:0] n13368_o;
  wire [76:0] n13369_o;
  wire [79:0] n13373_o;
  wire [63:0] n13375_o;
  wire n13385_o;
  wire [10:0] n13389_o;
  wire n13390_o;
  wire [10:0] n13392_o;
  wire n13393_o;
  wire [51:0] n13395_o;
  wire n13396_o;
  wire n13398_o;
  wire [10:0] n13399_o;
  wire [12:0] n13400_o;
  wire [12:0] n13402_o;
  wire n13403_o;
  wire [12:0] n13405_o;
  wire [9:0] n13407_o;
  wire [51:0] n13408_o;
  wire [61:0] n13409_o;
  wire [63:0] n13411_o;
  wire [1:0] n13412_o;
  wire [2:0] n13413_o;
  wire n13416_o;
  wire n13419_o;
  wire n13422_o;
  wire n13425_o;
  wire n13428_o;
  wire [4:0] n13430_o;
  reg [1:0] n13431_o;
  wire n13433_o;
  wire n13434_o;
  wire n13435_o;
  wire [1:0] n13438_o;
  wire [76:0] n13439_o;
  wire [76:0] n13440_o;
  wire [1:0] n13441_o;
  wire [76:0] n13442_o;
  wire [79:0] n13446_o;
  wire [12:0] n13448_o;
  wire [12:0] n13449_o;
  wire n13450_o;
  wire n13452_o;
  wire [12:0] n13454_o;
  wire [12:0] n13455_o;
  wire [12:0] n13456_o;
  wire [12:0] n13458_o;
  wire [12:0] n13459_o;
  wire n13460_o;
  wire n13462_o;
  wire [115:0] n13463_o;
  wire [239:0] n13464_o;
  wire [11:0] n13465_o;
  wire [115:0] n13466_o;
  wire [115:0] n13467_o;
  wire [239:0] n13468_o;
  wire [239:0] n13469_o;
  wire n13470_o;
  wire n13471_o;
  wire [7:0] n13472_o;
  wire [7:0] n13473_o;
  wire [11:0] n13474_o;
  wire [11:0] n13475_o;
  wire [1:0] n13476_o;
  wire [1:0] n13477_o;
  wire n13478_o;
  wire n13479_o;
  wire [31:0] n13483_o;
  wire [3:0] n13487_o;
  wire n13497_o;
  wire [24:0] n13499_o;
  wire n13500_o;
  wire [28:0] n13501_o;
  wire n13502_o;
  wire [55:0] n13503_o;
  wire n13504_o;
  wire n13505_o;
  wire n13506_o;
  wire n13507_o;
  wire n13508_o;
  wire [12:0] n13511_o;
  wire n13512_o;
  wire n13513_o;
  wire [12:0] n13516_o;
  wire [12:0] n13518_o;
  wire [12:0] n13520_o;
  wire [12:0] n13523_o;
  wire [12:0] n13524_o;
  wire [12:0] n13525_o;
  wire [12:0] n13526_o;
  wire n13527_o;
  wire n13530_o;
  wire n13532_o;
  wire n13535_o;
  wire [53:0] n13537_o;
  wire n13538_o;
  wire [55:0] n13539_o;
  wire [55:0] n13540_o;
  wire n13541_o;
  wire n13544_o;
  wire [55:0] n13546_o;
  wire [55:0] n13547_o;
  wire n13548_o;
  wire n13551_o;
  wire [1:0] n13556_o;
  wire [4:0] n13558_o;
  wire [264:0] n13560_o;
  wire [1:0] n13562_o;
  wire [4:0] n13564_o;
  wire [6:0] n13567_o;
  wire n13573_o;
  wire [4:0] n13574_o;
  wire n13575_o;
  wire n13576_o;
  wire n13577_o;
  wire [6:0] n13580_o;
  wire n13581_o;
  wire [6:0] n13585_o;
  wire [1:0] n13586_o;
  wire [6:0] n13587_o;
  wire [1:0] n13588_o;
  wire n13590_o;
  wire n13591_o;
  wire n13592_o;
  wire n13593_o;
  wire n13594_o;
  wire [6:0] n13597_o;
  wire [6:0] n13599_o;
  wire n13601_o;
  wire n13602_o;
  wire n13603_o;
  wire [6:0] n13606_o;
  wire n13608_o;
  wire [1:0] n13610_o;
  wire n13612_o;
  wire [6:0] n13615_o;
  wire n13617_o;
  wire n13621_o;
  wire [6:0] n13625_o;
  wire n13627_o;
  wire n13632_o;
  wire [721:0] n13634_o;
  wire n13635_o;
  wire n13636_o;
  wire [721:0] n13637_o;
  wire n13638_o;
  wire n13639_o;
  wire [1:0] n13641_o;
  wire n13644_o;
  wire n13648_o;
  wire n13650_o;
  wire n13651_o;
  wire n13656_o;
  wire n13659_o;
  wire n13663_o;
  wire [9:0] n13666_o;
  wire [9:0] n13667_o;
  wire [9:0] n13668_o;
  wire n13669_o;
  wire n13670_o;
  wire n13671_o;
  wire [721:0] n13672_o;
  wire n13673_o;
  wire n13674_o;
  wire [9:0] n13675_o;
  wire [9:0] n13676_o;
  wire [9:0] n13677_o;
  wire n13678_o;
  wire n13679_o;
  wire n13680_o;
  wire [721:0] n13681_o;
  wire n13682_o;
  wire n13683_o;
  wire [1:0] n13685_o;
  wire n13688_o;
  wire n13693_o;
  wire [721:0] n13694_o;
  wire n13695_o;
  wire n13696_o;
  wire [721:0] n13698_o;
  wire n13699_o;
  wire n13700_o;
  wire [1:0] n13703_o;
  wire [1:0] n13704_o;
  wire n13707_o;
  wire n13709_o;
  wire n13710_o;
  wire n13712_o;
  wire n13713_o;
  wire n13715_o;
  wire n13716_o;
  wire [14:0] n13717_o;
  reg [6:0] n13718_o;
  wire [2:0] n13719_o;
  wire [2:0] n13720_o;
  wire [2:0] n13721_o;
  reg [2:0] n13722_o;
  wire n13723_o;
  wire n13724_o;
  wire n13725_o;
  reg n13726_o;
  wire n13727_o;
  wire n13728_o;
  wire n13729_o;
  reg n13730_o;
  reg [1:0] n13731_o;
  reg n13734_o;
  wire [1:0] n13735_o;
  wire [6:0] n13736_o;
  wire [2:0] n13737_o;
  wire [2:0] n13738_o;
  wire [2:0] n13739_o;
  wire [2:0] n13740_o;
  wire [1:0] n13741_o;
  wire [1:0] n13742_o;
  wire [1:0] n13743_o;
  wire [1:0] n13744_o;
  wire [1:0] n13745_o;
  wire n13747_o;
  wire [4:0] n13749_o;
  wire n13751_o;
  wire [31:0] n13753_o;
  wire [2:0] n13758_o;
  wire [30:0] n13759_o;
  wire [31:0] n13760_o;
  wire n13762_o;
  wire [3:0] n13763_o;
  wire [3:0] n13765_o;
  wire [3:0] n13767_o;
  wire n13771_o;
  wire [3:0] n13772_o;
  wire [3:0] n13774_o;
  wire [3:0] n13776_o;
  wire n13780_o;
  wire [3:0] n13781_o;
  wire [3:0] n13783_o;
  wire [3:0] n13785_o;
  wire n13789_o;
  wire [3:0] n13790_o;
  wire [3:0] n13792_o;
  wire [3:0] n13794_o;
  wire n13798_o;
  wire [3:0] n13799_o;
  wire [3:0] n13801_o;
  wire [3:0] n13803_o;
  wire n13807_o;
  wire [3:0] n13808_o;
  wire [3:0] n13810_o;
  wire [3:0] n13812_o;
  wire n13816_o;
  wire [3:0] n13817_o;
  wire [3:0] n13819_o;
  wire [3:0] n13821_o;
  wire n13825_o;
  wire [3:0] n13826_o;
  wire [3:0] n13828_o;
  wire [3:0] n13830_o;
  wire [31:0] n13833_o;
  wire [31:0] n13835_o;
  wire [31:0] n13836_o;
  wire [31:0] n13837_o;
  wire n13841_o;
  localparam [3:0] n13844_o = 4'b0000;
  wire [79:0] n13845_o;
  wire [1:0] n13846_o;
  wire n13848_o;
  wire [79:0] n13849_o;
  wire [1:0] n13850_o;
  wire n13852_o;
  wire n13853_o;
  wire [79:0] n13854_o;
  wire [1:0] n13855_o;
  wire n13857_o;
  wire n13858_o;
  wire [79:0] n13859_o;
  wire [1:0] n13860_o;
  wire n13862_o;
  wire n13863_o;
  wire n13864_o;
  wire n13865_o;
  wire n13866_o;
  wire n13868_o;
  wire n13869_o;
  wire n13870_o;
  wire [79:0] n13872_o;
  wire [1:0] n13873_o;
  wire n13875_o;
  wire [79:0] n13876_o;
  wire [1:0] n13877_o;
  wire n13879_o;
  wire n13880_o;
  wire [79:0] n13881_o;
  wire [1:0] n13882_o;
  wire n13884_o;
  wire n13885_o;
  wire [79:0] n13886_o;
  wire [1:0] n13887_o;
  wire n13889_o;
  wire n13890_o;
  wire [79:0] n13891_o;
  wire [1:0] n13892_o;
  wire n13894_o;
  wire n13895_o;
  wire [79:0] n13896_o;
  wire [1:0] n13897_o;
  wire n13899_o;
  wire [79:0] n13900_o;
  wire [12:0] n13901_o;
  wire n13903_o;
  wire n13904_o;
  wire n13905_o;
  wire [6:0] n13911_o;
  wire n13912_o;
  wire n13913_o;
  wire n13914_o;
  wire n13915_o;
  wire [1:0] n13916_o;
  wire n13917_o;
  wire n13919_o;
  localparam [3:0] n13922_o = 4'b0000;
  wire [79:0] n13923_o;
  wire [1:0] n13924_o;
  wire n13926_o;
  wire [79:0] n13927_o;
  wire [1:0] n13928_o;
  wire n13930_o;
  wire n13931_o;
  wire [79:0] n13932_o;
  wire [1:0] n13933_o;
  wire n13935_o;
  wire n13936_o;
  wire n13937_o;
  wire n13938_o;
  wire n13939_o;
  wire n13941_o;
  wire n13942_o;
  wire n13943_o;
  wire [79:0] n13945_o;
  wire [1:0] n13946_o;
  wire n13948_o;
  wire [79:0] n13949_o;
  wire [1:0] n13950_o;
  wire n13952_o;
  wire n13953_o;
  wire [79:0] n13954_o;
  wire [1:0] n13955_o;
  wire n13957_o;
  wire n13958_o;
  wire [79:0] n13959_o;
  wire n13960_o;
  wire n13961_o;
  wire [79:0] n13962_o;
  wire [12:0] n13963_o;
  wire n13965_o;
  wire n13966_o;
  wire n13968_o;
  wire n13969_o;
  wire n13970_o;
  wire n13972_o;
  wire [79:0] n13975_o;
  wire [12:0] n13976_o;
  wire [79:0] n13977_o;
  wire [1:0] n13978_o;
  wire n13980_o;
  wire n13981_o;
  wire n13982_o;
  wire n13983_o;
  wire [79:0] n13984_o;
  wire [1:0] n13985_o;
  wire n13987_o;
  wire n13988_o;
  wire n13989_o;
  wire n13990_o;
  wire n13991_o;
  wire n13993_o;
  wire n13994_o;
  wire n13995_o;
  wire n13996_o;
  wire n13998_o;
  wire n13999_o;
  wire [79:0] n14001_o;
  wire [1:0] n14002_o;
  wire n14004_o;
  wire [79:0] n14005_o;
  wire [1:0] n14006_o;
  wire n14008_o;
  wire n14009_o;
  wire n14010_o;
  wire n14012_o;
  wire n14013_o;
  wire n14016_o;
  wire [79:0] n14018_o;
  wire [1:0] n14019_o;
  wire n14021_o;
  wire [79:0] n14022_o;
  wire [1:0] n14023_o;
  wire n14025_o;
  wire n14026_o;
  wire [79:0] n14028_o;
  wire n14029_o;
  wire [79:0] n14030_o;
  wire n14031_o;
  wire n14032_o;
  wire [79:0] n14033_o;
  wire n14034_o;
  wire [79:0] n14035_o;
  wire n14036_o;
  wire [1:0] n14037_o;
  wire [3:0] n14039_o;
  wire [79:0] n14040_o;
  wire [1:0] n14041_o;
  wire n14043_o;
  wire [79:0] n14044_o;
  wire n14045_o;
  wire n14046_o;
  wire [79:0] n14047_o;
  wire n14048_o;
  wire [1:0] n14049_o;
  wire [3:0] n14051_o;
  wire [79:0] n14052_o;
  wire [1:0] n14053_o;
  wire n14055_o;
  wire [79:0] n14056_o;
  wire [1:0] n14057_o;
  wire n14059_o;
  wire [79:0] n14061_o;
  wire n14062_o;
  wire [79:0] n14063_o;
  wire n14064_o;
  wire n14065_o;
  wire [1:0] n14066_o;
  wire [3:0] n14068_o;
  wire [3:0] n14069_o;
  wire [79:0] n14070_o;
  wire [1:0] n14071_o;
  wire n14073_o;
  wire [79:0] n14074_o;
  wire n14075_o;
  wire [79:0] n14076_o;
  wire n14077_o;
  wire n14078_o;
  wire [1:0] n14079_o;
  wire [3:0] n14081_o;
  wire [79:0] n14082_o;
  wire [1:0] n14083_o;
  wire n14085_o;
  wire [79:0] n14086_o;
  wire n14087_o;
  wire n14088_o;
  wire [79:0] n14089_o;
  wire n14090_o;
  wire [1:0] n14091_o;
  wire [3:0] n14093_o;
  wire n14094_o;
  wire [79:0] n14095_o;
  wire n14096_o;
  wire [79:0] n14097_o;
  wire n14098_o;
  wire n14099_o;
  wire [1:0] n14100_o;
  wire [3:0] n14102_o;
  wire [79:0] n14103_o;
  wire [12:0] n14104_o;
  wire [79:0] n14105_o;
  wire [12:0] n14106_o;
  wire n14107_o;
  wire [79:0] n14108_o;
  wire n14109_o;
  wire n14110_o;
  wire [79:0] n14111_o;
  wire n14112_o;
  wire [1:0] n14113_o;
  wire [3:0] n14115_o;
  wire [6:0] n14120_o;
  wire n14121_o;
  wire [3:0] n14122_o;
  wire [1:0] n14123_o;
  wire [6:0] n14124_o;
  wire n14125_o;
  wire [3:0] n14126_o;
  wire [1:0] n14127_o;
  wire [6:0] n14128_o;
  wire n14129_o;
  wire [3:0] n14130_o;
  wire [1:0] n14131_o;
  wire [6:0] n14132_o;
  wire n14133_o;
  wire [3:0] n14134_o;
  wire [1:0] n14135_o;
  wire [6:0] n14136_o;
  wire n14137_o;
  wire [3:0] n14138_o;
  wire [1:0] n14139_o;
  wire [6:0] n14140_o;
  wire n14141_o;
  wire [3:0] n14142_o;
  wire [1:0] n14143_o;
  wire [6:0] n14144_o;
  wire n14145_o;
  wire [3:0] n14146_o;
  wire [1:0] n14147_o;
  wire [6:0] n14148_o;
  wire n14149_o;
  wire [3:0] n14150_o;
  wire [1:0] n14151_o;
  wire [6:0] n14152_o;
  wire n14153_o;
  wire n14155_o;
  wire [3:0] n14156_o;
  wire [1:0] n14157_o;
  wire n14159_o;
  wire [6:0] n14160_o;
  wire n14161_o;
  wire n14162_o;
  wire n14163_o;
  wire n14164_o;
  wire [3:0] n14165_o;
  wire [1:0] n14166_o;
  wire n14168_o;
  wire [18:0] n14169_o;
  wire [3:0] n14170_o;
  wire [6:0] n14171_o;
  wire [251:0] n14172_o;
  wire [721:0] n14173_o;
  wire [3:0] n14174_o;
  wire n14176_o;
  wire [31:0] n14178_o;
  wire [4:0] n14183_o;
  wire [30:0] n14184_o;
  wire [31:0] n14185_o;
  wire n14187_o;
  wire n14188_o;
  wire n14189_o;
  wire n14190_o;
  wire n14192_o;
  wire n14193_o;
  wire n14194_o;
  wire n14195_o;
  wire n14197_o;
  wire n14198_o;
  wire n14199_o;
  wire n14200_o;
  wire n14202_o;
  wire n14203_o;
  wire n14204_o;
  wire n14205_o;
  wire n14207_o;
  wire n14208_o;
  wire n14209_o;
  wire n14210_o;
  wire n14212_o;
  wire n14213_o;
  wire n14214_o;
  wire n14215_o;
  wire n14217_o;
  wire n14218_o;
  wire n14219_o;
  wire n14220_o;
  wire n14222_o;
  wire n14223_o;
  wire n14224_o;
  wire n14225_o;
  wire n14227_o;
  wire n14228_o;
  wire n14229_o;
  wire n14230_o;
  wire n14232_o;
  wire n14233_o;
  wire n14234_o;
  wire n14235_o;
  wire n14237_o;
  wire n14238_o;
  wire n14239_o;
  wire n14240_o;
  wire n14242_o;
  wire n14243_o;
  wire n14244_o;
  wire n14245_o;
  wire n14247_o;
  wire n14248_o;
  wire n14249_o;
  wire n14250_o;
  wire n14252_o;
  wire n14253_o;
  wire n14254_o;
  wire n14255_o;
  wire n14257_o;
  wire n14258_o;
  wire n14259_o;
  wire n14260_o;
  wire n14262_o;
  wire n14263_o;
  wire n14264_o;
  wire n14265_o;
  wire n14267_o;
  wire n14268_o;
  wire n14269_o;
  wire n14270_o;
  wire n14272_o;
  wire n14273_o;
  wire n14274_o;
  wire n14275_o;
  wire n14277_o;
  wire n14278_o;
  wire n14279_o;
  wire n14280_o;
  wire n14282_o;
  wire n14283_o;
  wire n14284_o;
  wire n14285_o;
  wire n14287_o;
  wire n14288_o;
  wire n14289_o;
  wire n14290_o;
  wire n14292_o;
  wire n14293_o;
  wire n14294_o;
  wire n14295_o;
  wire n14297_o;
  wire n14298_o;
  wire n14299_o;
  wire n14300_o;
  wire n14302_o;
  wire n14303_o;
  wire n14304_o;
  wire n14305_o;
  wire n14307_o;
  wire n14308_o;
  wire n14309_o;
  wire n14310_o;
  wire n14312_o;
  wire n14313_o;
  wire n14314_o;
  wire n14315_o;
  wire n14317_o;
  wire n14318_o;
  wire n14319_o;
  wire n14320_o;
  wire n14322_o;
  wire n14323_o;
  wire n14324_o;
  wire n14325_o;
  wire n14327_o;
  wire n14328_o;
  wire n14329_o;
  wire n14330_o;
  wire n14332_o;
  wire n14333_o;
  wire n14334_o;
  wire n14335_o;
  wire n14337_o;
  wire n14338_o;
  wire n14339_o;
  wire n14340_o;
  wire n14342_o;
  wire n14343_o;
  wire n14344_o;
  wire n14345_o;
  wire n14349_o;
  wire [31:0] n14351_o;
  wire [2:0] n14356_o;
  wire [30:0] n14357_o;
  wire [31:0] n14358_o;
  wire n14359_o;
  wire n14360_o;
  wire n14362_o;
  wire [31:0] n14364_o;
  wire [3:0] n14369_o;
  wire [3:0] n14370_o;
  wire [3:0] n14371_o;
  wire n14375_o;
  wire [31:0] n14377_o;
  wire [3:0] n14382_o;
  wire [3:0] n14383_o;
  wire [3:0] n14384_o;
  wire n14388_o;
  wire [31:0] n14390_o;
  wire [3:0] n14395_o;
  wire [3:0] n14396_o;
  wire [3:0] n14397_o;
  wire n14401_o;
  wire [31:0] n14403_o;
  wire [3:0] n14408_o;
  wire [3:0] n14409_o;
  wire [3:0] n14410_o;
  wire n14414_o;
  wire [31:0] n14416_o;
  wire [3:0] n14421_o;
  wire [3:0] n14422_o;
  wire [3:0] n14423_o;
  wire n14427_o;
  wire [31:0] n14429_o;
  wire [3:0] n14434_o;
  wire [3:0] n14435_o;
  wire [3:0] n14436_o;
  wire n14440_o;
  wire [31:0] n14442_o;
  wire [3:0] n14447_o;
  wire [3:0] n14448_o;
  wire [3:0] n14449_o;
  wire n14453_o;
  wire [31:0] n14455_o;
  wire [3:0] n14460_o;
  wire [3:0] n14461_o;
  wire [3:0] n14462_o;
  wire [31:0] n14465_o;
  wire [31:0] n14466_o;
  wire n14471_o;
  wire n14472_o;
  wire [2:0] n14474_o;
  wire [3:0] n14476_o;
  wire n14482_o;
  wire [4:0] n14485_o;
  wire n14487_o;
  wire n14490_o;
  wire n14492_o;
  wire n14494_o;
  wire n14495_o;
  wire [1:0] n14496_o;
  wire n14498_o;
  wire [1:0] n14499_o;
  wire n14501_o;
  wire n14503_o;
  wire [5:0] n14504_o;
  wire [1:0] n14505_o;
  reg [1:0] n14506_o;
  wire [4:0] n14507_o;
  reg [4:0] n14508_o;
  reg [31:0] n14514_o;
  reg n14517_o;
  wire n14521_o;
  wire n14522_o;
  wire n14523_o;
  wire [7:0] n14524_o;
  wire [7:0] n14526_o;
  wire [7:0] n14528_o;
  wire n14529_o;
  wire [3:0] n14530_o;
  wire [3:0] n14531_o;
  wire [3:0] n14532_o;
  wire n14533_o;
  wire [3:0] n14534_o;
  wire [3:0] n14535_o;
  wire [3:0] n14536_o;
  wire n14537_o;
  wire [3:0] n14538_o;
  wire [3:0] n14539_o;
  wire [3:0] n14540_o;
  wire n14541_o;
  wire [3:0] n14542_o;
  wire [3:0] n14543_o;
  wire [3:0] n14544_o;
  wire n14545_o;
  wire [3:0] n14546_o;
  wire [3:0] n14547_o;
  wire [3:0] n14548_o;
  wire n14549_o;
  wire [3:0] n14550_o;
  wire [3:0] n14551_o;
  wire [3:0] n14552_o;
  wire n14553_o;
  wire [3:0] n14554_o;
  wire [3:0] n14555_o;
  wire [3:0] n14556_o;
  wire n14557_o;
  wire [3:0] n14558_o;
  wire [3:0] n14559_o;
  wire [3:0] n14560_o;
  wire n14564_o;
  wire [79:0] n14565_o;
  wire [1:0] n14566_o;
  wire [79:0] n14567_o;
  wire [12:0] n14568_o;
  wire n14570_o;
  wire n14572_o;
  wire n14574_o;
  wire [79:0] n14575_o;
  wire n14576_o;
  wire n14577_o;
  wire [79:0] n14578_o;
  wire n14579_o;
  wire n14580_o;
  wire [79:0] n14581_o;
  wire n14582_o;
  wire n14583_o;
  wire n14584_o;
  wire n14585_o;
  wire n14586_o;
  wire n14591_o;
  wire [79:0] n14592_o;
  wire [1:0] n14593_o;
  wire [79:0] n14594_o;
  wire n14595_o;
  wire [79:0] n14596_o;
  wire [12:0] n14597_o;
  wire [79:0] n14600_o;
  wire [1:0] n14601_o;
  wire n14603_o;
  wire n14604_o;
  wire n14605_o;
  wire n14606_o;
  wire n14608_o;
  wire n14609_o;
  wire n14612_o;
  wire [79:0] n14613_o;
  wire [1:0] n14614_o;
  wire n14616_o;
  wire [79:0] n14617_o;
  wire [12:0] n14618_o;
  wire n14620_o;
  wire [79:0] n14621_o;
  wire [12:0] n14622_o;
  wire [12:0] n14624_o;
  wire [1:0] n14626_o;
  wire [2:0] n14628_o;
  wire [6:0] n14629_o;
  wire [12:0] n14630_o;
  wire [2:0] n14631_o;
  wire [2:0] n14632_o;
  wire [2:0] n14633_o;
  wire [2:0] n14634_o;
  wire n14637_o;
  wire [6:0] n14638_o;
  wire [12:0] n14639_o;
  wire [2:0] n14640_o;
  wire [2:0] n14641_o;
  wire [2:0] n14642_o;
  wire [2:0] n14643_o;
  wire n14645_o;
  wire n14647_o;
  wire [79:0] n14648_o;
  wire [1:0] n14649_o;
  wire [79:0] n14650_o;
  wire n14651_o;
  wire [79:0] n14652_o;
  wire [12:0] n14653_o;
  wire [79:0] n14656_o;
  wire [1:0] n14657_o;
  wire n14659_o;
  wire n14660_o;
  wire n14661_o;
  wire n14662_o;
  wire n14664_o;
  wire n14665_o;
  wire n14668_o;
  wire [79:0] n14669_o;
  wire [1:0] n14670_o;
  wire n14672_o;
  wire [79:0] n14673_o;
  wire [12:0] n14674_o;
  wire n14676_o;
  wire [79:0] n14677_o;
  wire [12:0] n14678_o;
  wire [12:0] n14680_o;
  wire [79:0] n14682_o;
  wire [12:0] n14683_o;
  wire n14685_o;
  wire [6:0] n14688_o;
  wire [6:0] n14689_o;
  wire [12:0] n14690_o;
  wire [6:0] n14691_o;
  wire n14692_o;
  wire n14695_o;
  wire n14697_o;
  wire [79:0] n14698_o;
  wire [1:0] n14699_o;
  wire [79:0] n14700_o;
  wire n14701_o;
  wire [79:0] n14702_o;
  wire [12:0] n14703_o;
  wire [79:0] n14706_o;
  wire [1:0] n14707_o;
  wire n14709_o;
  wire n14710_o;
  wire n14711_o;
  wire n14712_o;
  wire n14714_o;
  wire n14715_o;
  wire n14718_o;
  wire [79:0] n14720_o;
  wire [1:0] n14721_o;
  wire n14723_o;
  wire [79:0] n14724_o;
  wire [12:0] n14725_o;
  wire n14727_o;
  wire n14728_o;
  wire n14729_o;
  wire [79:0] n14730_o;
  wire [12:0] n14731_o;
  wire n14733_o;
  wire n14734_o;
  wire n14735_o;
  wire [79:0] n14737_o;
  wire [12:0] n14738_o;
  wire n14740_o;
  wire [79:0] n14741_o;
  wire [12:0] n14742_o;
  wire [12:0] n14744_o;
  wire n14745_o;
  wire [79:0] n14746_o;
  wire n14747_o;
  wire n14748_o;
  wire [6:0] n14751_o;
  wire [79:0] n14752_o;
  wire [12:0] n14753_o;
  wire [12:0] n14755_o;
  wire [6:0] n14757_o;
  wire [12:0] n14758_o;
  wire [6:0] n14759_o;
  wire [12:0] n14760_o;
  wire n14762_o;
  wire n14765_o;
  wire n14767_o;
  wire n14768_o;
  wire [2:0] n14769_o;
  reg [6:0] n14771_o;
  reg [12:0] n14773_o;
  reg n14777_o;
  wire n14779_o;
  wire n14781_o;
  wire n14782_o;
  wire [79:0] n14783_o;
  wire n14784_o;
  wire n14785_o;
  wire n14789_o;
  wire n14792_o;
  wire n14793_o;
  wire [79:0] n14794_o;
  wire [1:0] n14795_o;
  wire [79:0] n14799_o;
  wire [1:0] n14800_o;
  wire n14802_o;
  wire [6:0] n14804_o;
  wire n14807_o;
  wire n14809_o;
  wire [79:0] n14810_o;
  wire n14811_o;
  wire [79:0] n14812_o;
  wire [1:0] n14813_o;
  wire [79:0] n14814_o;
  wire [12:0] n14815_o;
  wire [79:0] n14820_o;
  wire n14821_o;
  wire [79:0] n14822_o;
  wire n14823_o;
  wire n14824_o;
  wire n14825_o;
  wire n14826_o;
  wire [79:0] n14827_o;
  wire [1:0] n14828_o;
  wire n14830_o;
  wire [79:0] n14831_o;
  wire [1:0] n14832_o;
  wire n14834_o;
  wire n14835_o;
  wire n14836_o;
  wire n14837_o;
  wire n14839_o;
  wire n14840_o;
  wire [79:0] n14841_o;
  wire [12:0] n14842_o;
  wire [79:0] n14843_o;
  wire [12:0] n14844_o;
  wire [12:0] n14845_o;
  wire [79:0] n14846_o;
  wire n14847_o;
  wire n14848_o;
  wire n14849_o;
  wire [79:0] n14850_o;
  wire [12:0] n14851_o;
  wire [79:0] n14852_o;
  wire [12:0] n14853_o;
  wire n14854_o;
  wire [6:0] n14858_o;
  wire n14859_o;
  wire [6:0] n14861_o;
  wire n14862_o;
  wire [12:0] n14863_o;
  wire n14864_o;
  wire [79:0] n14865_o;
  wire [1:0] n14866_o;
  wire n14868_o;
  wire [79:0] n14869_o;
  wire [1:0] n14870_o;
  wire n14872_o;
  wire n14873_o;
  wire [79:0] n14875_o;
  wire [1:0] n14876_o;
  wire n14878_o;
  wire [79:0] n14879_o;
  wire [1:0] n14880_o;
  wire n14882_o;
  wire n14883_o;
  wire n14884_o;
  wire n14885_o;
  wire [79:0] n14887_o;
  wire [1:0] n14888_o;
  wire n14890_o;
  wire [79:0] n14891_o;
  wire [1:0] n14892_o;
  wire n14894_o;
  wire n14895_o;
  wire n14896_o;
  wire n14897_o;
  wire n14898_o;
  wire n14899_o;
  wire n14900_o;
  wire [79:0] n14901_o;
  wire [1:0] n14902_o;
  wire n14904_o;
  wire [79:0] n14905_o;
  wire [1:0] n14906_o;
  wire n14908_o;
  wire n14909_o;
  wire n14913_o;
  wire n14914_o;
  wire [6:0] n14916_o;
  wire [1:0] n14917_o;
  wire n14918_o;
  wire n14919_o;
  wire [6:0] n14920_o;
  wire n14921_o;
  wire [1:0] n14922_o;
  wire n14923_o;
  wire n14924_o;
  wire n14927_o;
  wire [6:0] n14928_o;
  wire n14929_o;
  wire n14930_o;
  wire n14931_o;
  wire [1:0] n14932_o;
  wire n14933_o;
  wire n14934_o;
  wire n14936_o;
  wire n14939_o;
  wire [6:0] n14940_o;
  wire n14941_o;
  wire n14942_o;
  wire n14943_o;
  wire [1:0] n14944_o;
  wire n14945_o;
  wire n14946_o;
  wire n14948_o;
  wire n14950_o;
  wire [6:0] n14951_o;
  wire n14952_o;
  wire n14953_o;
  wire n14954_o;
  wire n14955_o;
  wire n14956_o;
  wire n14957_o;
  wire n14958_o;
  wire n14959_o;
  wire n14960_o;
  wire n14961_o;
  wire n14962_o;
  wire n14963_o;
  wire [1:0] n14964_o;
  wire n14965_o;
  wire n14966_o;
  wire n14967_o;
  wire n14969_o;
  wire n14971_o;
  wire n14973_o;
  wire [79:0] n14974_o;
  wire n14975_o;
  wire [79:0] n14976_o;
  wire n14977_o;
  wire n14978_o;
  wire [79:0] n14979_o;
  wire [1:0] n14980_o;
  wire [79:0] n14985_o;
  wire [1:0] n14986_o;
  wire n14988_o;
  wire [79:0] n14989_o;
  wire [1:0] n14990_o;
  wire n14992_o;
  wire n14993_o;
  wire [79:0] n14994_o;
  wire [12:0] n14995_o;
  wire [79:0] n14996_o;
  wire [12:0] n14997_o;
  wire [12:0] n14998_o;
  wire n14999_o;
  wire n15000_o;
  wire n15002_o;
  wire n15003_o;
  wire n15007_o;
  wire [6:0] n15008_o;
  wire n15009_o;
  wire [6:0] n15010_o;
  wire [79:0] n15011_o;
  wire [1:0] n15012_o;
  wire n15014_o;
  wire [79:0] n15015_o;
  wire [1:0] n15016_o;
  wire n15018_o;
  wire n15019_o;
  wire [79:0] n15021_o;
  wire [1:0] n15022_o;
  wire n15024_o;
  wire [79:0] n15025_o;
  wire [1:0] n15026_o;
  wire n15028_o;
  wire n15029_o;
  wire [79:0] n15030_o;
  wire [1:0] n15031_o;
  wire n15033_o;
  wire [79:0] n15034_o;
  wire [1:0] n15035_o;
  wire n15037_o;
  wire n15038_o;
  wire n15039_o;
  wire [79:0] n15041_o;
  wire [1:0] n15042_o;
  wire n15044_o;
  wire [79:0] n15045_o;
  wire [1:0] n15046_o;
  wire n15048_o;
  wire n15049_o;
  wire [79:0] n15051_o;
  wire n15052_o;
  wire [6:0] n15054_o;
  wire [1:0] n15055_o;
  wire n15056_o;
  wire n15057_o;
  wire n15060_o;
  wire [6:0] n15061_o;
  wire n15062_o;
  wire n15063_o;
  wire [1:0] n15064_o;
  wire n15065_o;
  wire n15066_o;
  wire n15068_o;
  wire n15071_o;
  wire [6:0] n15072_o;
  wire n15073_o;
  wire n15074_o;
  wire [1:0] n15075_o;
  wire n15076_o;
  wire n15077_o;
  wire n15079_o;
  wire n15081_o;
  wire n15082_o;
  wire [6:0] n15083_o;
  wire n15084_o;
  wire n15085_o;
  wire [12:0] n15086_o;
  wire [12:0] n15087_o;
  wire [1:0] n15088_o;
  wire n15089_o;
  wire n15090_o;
  wire n15092_o;
  wire n15094_o;
  wire n15096_o;
  wire [79:0] n15097_o;
  wire [1:0] n15098_o;
  wire [79:0] n15103_o;
  wire n15104_o;
  wire [79:0] n15105_o;
  wire n15106_o;
  wire n15107_o;
  wire [79:0] n15108_o;
  wire [12:0] n15109_o;
  wire [79:0] n15110_o;
  wire [12:0] n15111_o;
  wire [12:0] n15112_o;
  wire [79:0] n15114_o;
  wire [1:0] n15115_o;
  wire n15117_o;
  wire [79:0] n15118_o;
  wire [1:0] n15119_o;
  wire n15121_o;
  wire n15122_o;
  wire n15123_o;
  wire n15124_o;
  wire n15126_o;
  wire n15127_o;
  wire [6:0] n15131_o;
  wire n15132_o;
  wire [6:0] n15133_o;
  wire n15134_o;
  wire [79:0] n15135_o;
  wire [1:0] n15136_o;
  wire n15138_o;
  wire [79:0] n15139_o;
  wire [1:0] n15140_o;
  wire n15142_o;
  wire n15143_o;
  wire [79:0] n15145_o;
  wire [1:0] n15146_o;
  wire n15148_o;
  wire [79:0] n15149_o;
  wire [1:0] n15150_o;
  wire n15152_o;
  wire n15155_o;
  wire n15156_o;
  wire [1:0] n15157_o;
  wire n15160_o;
  wire [79:0] n15161_o;
  wire [1:0] n15162_o;
  wire n15164_o;
  wire [79:0] n15165_o;
  wire [1:0] n15166_o;
  wire n15168_o;
  wire [79:0] n15170_o;
  wire [1:0] n15171_o;
  wire n15173_o;
  wire n15176_o;
  wire n15178_o;
  wire n15179_o;
  wire [1:0] n15180_o;
  wire n15182_o;
  wire n15185_o;
  wire n15187_o;
  wire [1:0] n15188_o;
  wire n15190_o;
  wire n15192_o;
  wire n15193_o;
  wire n15194_o;
  wire n15196_o;
  wire [1:0] n15197_o;
  wire n15199_o;
  wire n15200_o;
  wire [1:0] n15201_o;
  wire [6:0] n15202_o;
  wire [1:0] n15203_o;
  wire [1:0] n15204_o;
  wire [1:0] n15205_o;
  wire n15208_o;
  wire n15210_o;
  wire n15212_o;
  wire [6:0] n15213_o;
  wire [1:0] n15214_o;
  wire [1:0] n15215_o;
  wire [1:0] n15216_o;
  wire n15217_o;
  wire n15219_o;
  wire n15221_o;
  wire n15223_o;
  wire n15225_o;
  wire [79:0] n15228_o;
  wire [1:0] n15229_o;
  wire n15231_o;
  wire [79:0] n15232_o;
  wire n15233_o;
  wire n15234_o;
  wire [79:0] n15235_o;
  wire [1:0] n15236_o;
  wire n15238_o;
  wire n15239_o;
  wire n15240_o;
  wire [1:0] n15243_o;
  wire n15247_o;
  wire [79:0] n15248_o;
  wire [1:0] n15249_o;
  wire [79:0] n15250_o;
  wire n15251_o;
  wire [79:0] n15255_o;
  wire [1:0] n15256_o;
  wire [79:0] n15257_o;
  wire [12:0] n15258_o;
  wire [79:0] n15259_o;
  wire n15260_o;
  wire n15262_o;
  wire n15263_o;
  wire n15265_o;
  wire n15266_o;
  wire [6:0] n15270_o;
  wire [12:0] n15271_o;
  wire [6:0] n15272_o;
  wire [12:0] n15273_o;
  wire [6:0] n15274_o;
  wire n15275_o;
  wire n15276_o;
  wire [12:0] n15277_o;
  wire n15280_o;
  wire n15282_o;
  wire n15285_o;
  wire n15287_o;
  wire [79:0] n15288_o;
  wire n15289_o;
  wire n15291_o;
  wire n15292_o;
  wire n15295_o;
  wire n15297_o;
  wire [3:0] n15298_o;
  reg [6:0] n15300_o;
  wire n15301_o;
  reg n15303_o;
  wire [12:0] n15304_o;
  reg [12:0] n15306_o;
  reg [12:0] n15308_o;
  reg n15313_o;
  reg n15316_o;
  wire n15318_o;
  wire [79:0] n15319_o;
  wire [1:0] n15320_o;
  wire [79:0] n15321_o;
  wire n15322_o;
  wire [79:0] n15326_o;
  wire [1:0] n15327_o;
  wire [79:0] n15328_o;
  wire [12:0] n15329_o;
  wire [12:0] n15330_o;
  wire n15331_o;
  wire n15332_o;
  wire [6:0] n15335_o;
  wire n15337_o;
  wire n15340_o;
  wire n15343_o;
  wire n15346_o;
  wire [3:0] n15347_o;
  reg [6:0] n15349_o;
  reg [1:0] n15351_o;
  wire [12:0] n15352_o;
  reg [12:0] n15354_o;
  reg n15359_o;
  reg n15363_o;
  wire n15365_o;
  wire [79:0] n15366_o;
  wire [1:0] n15367_o;
  wire [79:0] n15368_o;
  wire n15369_o;
  wire [79:0] n15374_o;
  wire [1:0] n15375_o;
  wire [79:0] n15376_o;
  wire [12:0] n15377_o;
  wire [79:0] n15378_o;
  wire n15379_o;
  wire n15381_o;
  wire n15382_o;
  wire n15384_o;
  wire n15385_o;
  wire [6:0] n15388_o;
  wire [6:0] n15389_o;
  wire [6:0] n15390_o;
  wire n15391_o;
  wire n15392_o;
  wire n15395_o;
  wire n15397_o;
  wire n15400_o;
  wire [79:0] n15401_o;
  wire n15402_o;
  wire n15405_o;
  wire n15406_o;
  wire [1:0] n15407_o;
  wire n15410_o;
  wire n15412_o;
  wire n15415_o;
  wire [3:0] n15416_o;
  reg [6:0] n15418_o;
  wire n15419_o;
  reg n15421_o;
  reg [1:0] n15423_o;
  wire [12:0] n15424_o;
  reg [12:0] n15426_o;
  reg n15431_o;
  reg n15435_o;
  reg n15438_o;
  wire n15440_o;
  wire [79:0] n15441_o;
  wire n15442_o;
  wire [79:0] n15443_o;
  wire [1:0] n15444_o;
  wire [79:0] n15445_o;
  wire [12:0] n15446_o;
  wire [79:0] n15452_o;
  wire n15453_o;
  wire [79:0] n15454_o;
  wire n15455_o;
  wire n15456_o;
  wire [79:0] n15457_o;
  wire n15458_o;
  wire n15459_o;
  wire n15460_o;
  wire n15461_o;
  wire [79:0] n15462_o;
  wire [1:0] n15463_o;
  wire n15465_o;
  wire [79:0] n15466_o;
  wire [1:0] n15467_o;
  wire n15469_o;
  wire n15470_o;
  wire [79:0] n15471_o;
  wire [1:0] n15472_o;
  wire n15474_o;
  wire [79:0] n15475_o;
  wire [1:0] n15476_o;
  wire n15478_o;
  wire n15479_o;
  wire n15480_o;
  wire n15481_o;
  wire [79:0] n15482_o;
  wire [12:0] n15483_o;
  wire [79:0] n15484_o;
  wire [12:0] n15485_o;
  wire [12:0] n15486_o;
  wire n15487_o;
  wire n15488_o;
  wire n15490_o;
  wire n15491_o;
  wire [79:0] n15493_o;
  wire [1:0] n15494_o;
  wire n15496_o;
  wire [79:0] n15497_o;
  wire n15498_o;
  wire [79:0] n15499_o;
  wire n15500_o;
  wire n15501_o;
  wire n15502_o;
  wire n15503_o;
  wire n15507_o;
  wire n15508_o;
  wire [79:0] n15509_o;
  wire n15510_o;
  wire n15511_o;
  wire n15512_o;
  wire n15513_o;
  wire n15514_o;
  wire n15515_o;
  wire [79:0] n15518_o;
  wire [12:0] n15519_o;
  wire [12:0] n15520_o;
  wire [12:0] n15522_o;
  wire [79:0] n15523_o;
  wire n15524_o;
  wire [79:0] n15525_o;
  wire n15526_o;
  wire n15527_o;
  wire n15528_o;
  wire n15529_o;
  wire n15530_o;
  wire n15531_o;
  wire [79:0] n15532_o;
  wire [12:0] n15533_o;
  wire n15535_o;
  wire [25:0] n15536_o;
  wire [6:0] n15537_o;
  wire n15538_o;
  wire [25:0] n15539_o;
  wire [25:0] n15540_o;
  wire n15541_o;
  wire [6:0] n15542_o;
  wire n15543_o;
  wire [25:0] n15544_o;
  wire [25:0] n15545_o;
  wire n15546_o;
  wire n15547_o;
  wire n15548_o;
  wire n15549_o;
  wire n15550_o;
  wire [6:0] n15551_o;
  wire n15552_o;
  wire [25:0] n15553_o;
  wire [25:0] n15554_o;
  wire n15555_o;
  wire n15556_o;
  wire n15557_o;
  wire n15558_o;
  wire n15559_o;
  wire [6:0] n15560_o;
  wire n15561_o;
  wire [25:0] n15562_o;
  wire [25:0] n15563_o;
  wire n15564_o;
  wire n15565_o;
  wire n15566_o;
  wire n15567_o;
  wire [79:0] n15568_o;
  wire [1:0] n15569_o;
  wire n15571_o;
  wire [79:0] n15572_o;
  wire [1:0] n15573_o;
  wire n15575_o;
  wire n15576_o;
  wire [79:0] n15577_o;
  wire [1:0] n15578_o;
  wire n15580_o;
  wire n15581_o;
  wire [79:0] n15583_o;
  wire [1:0] n15584_o;
  wire n15586_o;
  wire [79:0] n15587_o;
  wire [1:0] n15588_o;
  wire n15590_o;
  wire n15591_o;
  wire [79:0] n15592_o;
  wire [1:0] n15593_o;
  wire n15595_o;
  wire [79:0] n15596_o;
  wire [1:0] n15597_o;
  wire n15599_o;
  wire n15600_o;
  wire n15601_o;
  wire [79:0] n15603_o;
  wire [1:0] n15604_o;
  wire n15606_o;
  wire [79:0] n15607_o;
  wire [1:0] n15608_o;
  wire n15610_o;
  wire n15611_o;
  wire [79:0] n15612_o;
  wire [1:0] n15613_o;
  wire n15615_o;
  wire n15616_o;
  wire n15617_o;
  wire [79:0] n15620_o;
  wire n15621_o;
  wire [79:0] n15622_o;
  wire n15623_o;
  wire n15624_o;
  wire n15625_o;
  wire n15626_o;
  wire [2:0] n15627_o;
  wire n15628_o;
  wire n15629_o;
  wire [2:0] n15630_o;
  wire [2:0] n15631_o;
  wire n15634_o;
  wire n15637_o;
  wire [79:0] n15639_o;
  wire [1:0] n15640_o;
  wire n15642_o;
  wire n15643_o;
  wire n15644_o;
  wire n15645_o;
  wire n15646_o;
  wire n15647_o;
  wire [79:0] n15648_o;
  wire n15649_o;
  wire n15650_o;
  wire n15651_o;
  wire n15652_o;
  wire n15653_o;
  wire n15654_o;
  wire n15655_o;
  wire n15656_o;
  wire [6:0] n15658_o;
  wire n15660_o;
  wire [2:0] n15661_o;
  wire [2:0] n15662_o;
  wire [1:0] n15663_o;
  wire n15664_o;
  wire n15665_o;
  wire n15667_o;
  wire n15669_o;
  wire [6:0] n15670_o;
  wire n15671_o;
  wire n15672_o;
  wire n15673_o;
  wire n15674_o;
  wire [2:0] n15675_o;
  wire [2:0] n15676_o;
  wire [1:0] n15677_o;
  wire n15678_o;
  wire n15679_o;
  wire n15681_o;
  wire n15683_o;
  wire [6:0] n15684_o;
  wire n15685_o;
  wire n15686_o;
  wire n15687_o;
  wire n15688_o;
  wire [2:0] n15689_o;
  wire [2:0] n15690_o;
  wire [1:0] n15691_o;
  wire n15692_o;
  wire n15693_o;
  wire n15695_o;
  wire n15697_o;
  wire n15698_o;
  wire [6:0] n15699_o;
  wire n15700_o;
  wire n15701_o;
  wire n15702_o;
  wire n15703_o;
  wire n15704_o;
  wire n15705_o;
  wire [1:0] n15706_o;
  wire [1:0] n15707_o;
  wire [25:0] n15708_o;
  wire [25:0] n15709_o;
  wire n15710_o;
  wire n15711_o;
  wire n15712_o;
  wire n15713_o;
  wire n15714_o;
  wire n15715_o;
  wire n15716_o;
  wire n15717_o;
  wire [1:0] n15718_o;
  wire n15719_o;
  wire n15720_o;
  wire n15722_o;
  wire n15724_o;
  wire n15727_o;
  wire n15729_o;
  wire [1:0] n15732_o;
  wire n15734_o;
  wire n15735_o;
  wire n15736_o;
  wire n15737_o;
  wire n15738_o;
  wire [79:0] n15739_o;
  wire [1:0] n15740_o;
  wire n15742_o;
  wire n15743_o;
  wire [12:0] n15748_o;
  wire [79:0] n15749_o;
  wire [12:0] n15750_o;
  wire n15751_o;
  wire n15753_o;
  wire [6:0] n15756_o;
  wire n15757_o;
  wire n15758_o;
  wire n15759_o;
  wire n15760_o;
  wire n15761_o;
  wire [1:0] n15762_o;
  wire [6:0] n15764_o;
  wire n15765_o;
  wire n15766_o;
  wire n15767_o;
  wire n15768_o;
  wire n15769_o;
  wire [1:0] n15770_o;
  wire n15771_o;
  wire [6:0] n15775_o;
  wire n15776_o;
  wire [6:0] n15777_o;
  wire n15778_o;
  wire n15779_o;
  wire n15780_o;
  wire n15781_o;
  wire n15782_o;
  wire n15783_o;
  wire n15785_o;
  wire n15786_o;
  wire n15789_o;
  wire n15790_o;
  wire n15791_o;
  wire [12:0] n15792_o;
  wire [12:0] n15793_o;
  wire [12:0] n15794_o;
  wire [12:0] n15795_o;
  wire n15799_o;
  wire n15802_o;
  wire n15803_o;
  wire n15804_o;
  wire [79:0] n15805_o;
  wire [1:0] n15806_o;
  wire n15808_o;
  wire n15809_o;
  wire [12:0] n15814_o;
  wire [79:0] n15815_o;
  wire [12:0] n15816_o;
  wire n15817_o;
  wire n15819_o;
  wire [6:0] n15822_o;
  wire n15823_o;
  wire n15824_o;
  wire n15825_o;
  wire n15826_o;
  wire n15827_o;
  wire [1:0] n15828_o;
  wire n15830_o;
  wire [79:0] n15831_o;
  wire [12:0] n15832_o;
  wire [79:0] n15833_o;
  wire [12:0] n15834_o;
  wire [12:0] n15835_o;
  wire [79:0] n15836_o;
  wire [12:0] n15837_o;
  wire n15841_o;
  wire n15842_o;
  wire n15843_o;
  wire [1:0] n15846_o;
  wire n15849_o;
  wire n15850_o;
  wire n15851_o;
  wire n15852_o;
  wire n15853_o;
  wire n15854_o;
  wire n15858_o;
  wire n15859_o;
  wire n15860_o;
  wire n15861_o;
  wire n15863_o;
  wire [6:0] n15866_o;
  wire n15867_o;
  wire n15869_o;
  wire n15870_o;
  wire n15871_o;
  wire n15872_o;
  wire n15873_o;
  wire n15874_o;
  wire n15876_o;
  wire n15877_o;
  wire n15878_o;
  wire n15879_o;
  wire n15880_o;
  wire n15881_o;
  wire [2:0] n15883_o;
  wire [6:0] n15884_o;
  wire [2:0] n15885_o;
  wire [2:0] n15886_o;
  wire n15889_o;
  wire n15892_o;
  wire [6:0] n15893_o;
  wire [2:0] n15894_o;
  wire [2:0] n15895_o;
  wire n15897_o;
  wire n15899_o;
  wire n15902_o;
  wire [1:0] n15905_o;
  wire [6:0] n15906_o;
  wire [2:0] n15907_o;
  wire [2:0] n15908_o;
  wire n15910_o;
  wire n15912_o;
  wire n15914_o;
  wire [1:0] n15916_o;
  wire n15919_o;
  wire n15922_o;
  wire [6:0] n15923_o;
  wire n15924_o;
  wire n15925_o;
  wire [1:0] n15926_o;
  wire [1:0] n15927_o;
  wire [1:0] n15928_o;
  wire n15930_o;
  wire n15932_o;
  wire n15934_o;
  wire n15936_o;
  wire n15939_o;
  wire n15940_o;
  wire [79:0] n15941_o;
  wire n15942_o;
  wire n15943_o;
  wire [79:0] n15944_o;
  wire n15945_o;
  wire [1:0] n15946_o;
  wire [3:0] n15948_o;
  wire n15949_o;
  wire n15950_o;
  wire [79:0] n15952_o;
  wire n15953_o;
  wire [79:0] n15954_o;
  wire n15955_o;
  wire n15956_o;
  wire [1:0] n15957_o;
  wire [3:0] n15959_o;
  wire [3:0] n15960_o;
  wire [3:0] n15961_o;
  wire [721:0] n15962_o;
  wire [3:0] n15963_o;
  wire n15967_o;
  wire n15968_o;
  wire n15969_o;
  wire [6:0] n15971_o;
  wire n15973_o;
  wire [79:0] n15974_o;
  wire n15975_o;
  wire n15976_o;
  wire n15977_o;
  wire n15978_o;
  wire n15979_o;
  wire n15980_o;
  wire [12:0] n15981_o;
  wire [79:0] n15982_o;
  wire [12:0] n15983_o;
  wire [12:0] n15984_o;
  wire n15985_o;
  wire n15986_o;
  wire [6:0] n15989_o;
  wire n15990_o;
  wire n15992_o;
  wire [12:0] n15993_o;
  wire [12:0] n15995_o;
  wire n15998_o;
  wire n16002_o;
  wire n16003_o;
  wire n16004_o;
  wire n16005_o;
  wire [6:0] n16007_o;
  wire n16009_o;
  wire n16010_o;
  wire n16011_o;
  wire n16012_o;
  wire n16013_o;
  wire n16014_o;
  wire n16015_o;
  wire [1:0] n16018_o;
  wire n16021_o;
  wire n16023_o;
  wire n16024_o;
  wire n16025_o;
  wire n16028_o;
  wire n16032_o;
  wire n16033_o;
  wire n16034_o;
  wire n16035_o;
  wire n16036_o;
  wire n16037_o;
  wire n16038_o;
  wire n16039_o;
  wire n16040_o;
  wire n16041_o;
  wire n16043_o;
  wire n16044_o;
  wire n16045_o;
  wire [1:0] n16048_o;
  wire [2:0] n16049_o;
  wire [2:0] n16050_o;
  wire [2:0] n16051_o;
  wire n16054_o;
  wire n16057_o;
  wire [2:0] n16058_o;
  wire n16060_o;
  wire [6:0] n16063_o;
  wire n16066_o;
  wire [1:0] n16068_o;
  wire [6:0] n16069_o;
  wire n16071_o;
  wire n16073_o;
  wire n16075_o;
  wire n16077_o;
  wire n16079_o;
  wire n16081_o;
  wire n16082_o;
  wire n16083_o;
  wire n16084_o;
  wire [6:0] n16087_o;
  wire n16088_o;
  wire n16089_o;
  wire [6:0] n16092_o;
  wire [6:0] n16093_o;
  wire n16095_o;
  wire [1:0] n16096_o;
  wire n16098_o;
  wire [1:0] n16101_o;
  wire n16102_o;
  wire n16103_o;
  wire n16104_o;
  wire [1:0] n16106_o;
  wire [1:0] n16108_o;
  wire [2:0] n16110_o;
  wire [6:0] n16111_o;
  wire [2:0] n16112_o;
  wire [2:0] n16113_o;
  wire n16115_o;
  wire n16116_o;
  wire n16117_o;
  wire [1:0] n16119_o;
  wire n16121_o;
  wire [6:0] n16124_o;
  wire [6:0] n16125_o;
  wire n16126_o;
  wire n16128_o;
  wire n16129_o;
  wire n16130_o;
  wire n16131_o;
  wire [1:0] n16136_o;
  wire [6:0] n16137_o;
  wire n16138_o;
  wire n16140_o;
  wire n16141_o;
  wire n16142_o;
  wire [6:0] n16144_o;
  wire n16146_o;
  wire n16147_o;
  wire n16148_o;
  wire n16149_o;
  wire n16152_o;
  wire n16153_o;
  wire n16156_o;
  wire n16160_o;
  wire n16161_o;
  wire n16162_o;
  wire [79:0] n16163_o;
  wire [1:0] n16164_o;
  wire n16166_o;
  wire n16167_o;
  wire n16168_o;
  wire n16169_o;
  wire n16170_o;
  wire [79:0] n16173_o;
  wire [12:0] n16174_o;
  wire [6:0] n16176_o;
  wire n16177_o;
  wire [12:0] n16178_o;
  wire [1:0] n16179_o;
  wire n16181_o;
  wire n16182_o;
  wire [11:0] n16183_o;
  wire [12:0] n16184_o;
  wire [12:0] n16185_o;
  wire n16189_o;
  wire n16195_o;
  wire n16199_o;
  wire n16200_o;
  wire n16201_o;
  wire [1:0] n16206_o;
  wire [6:0] n16207_o;
  wire n16208_o;
  wire n16210_o;
  wire n16211_o;
  wire n16212_o;
  wire [6:0] n16214_o;
  wire n16216_o;
  wire n16221_o;
  wire n16222_o;
  wire n16223_o;
  wire [6:0] n16226_o;
  wire n16227_o;
  wire n16229_o;
  wire n16230_o;
  wire n16231_o;
  wire [1:0] n16233_o;
  wire [1:0] n16235_o;
  wire [1:0] n16236_o;
  wire n16238_o;
  wire [6:0] n16242_o;
  wire n16243_o;
  wire [1:0] n16246_o;
  wire [2:0] n16247_o;
  wire [6:0] n16248_o;
  wire [2:0] n16249_o;
  wire [2:0] n16250_o;
  wire n16252_o;
  wire n16253_o;
  wire n16254_o;
  wire [6:0] n16257_o;
  wire n16258_o;
  wire n16260_o;
  wire n16261_o;
  wire n16262_o;
  wire [6:0] n16264_o;
  wire n16266_o;
  wire n16267_o;
  wire [11:0] n16268_o;
  wire [12:0] n16269_o;
  wire n16274_o;
  wire n16275_o;
  wire n16276_o;
  wire n16277_o;
  wire [6:0] n16279_o;
  wire n16281_o;
  wire n16282_o;
  wire n16283_o;
  wire n16284_o;
  wire n16287_o;
  wire n16288_o;
  wire n16291_o;
  wire n16295_o;
  wire [63:0] n16297_o;
  wire n16298_o;
  wire [2:0] n16299_o;
  wire n16300_o;
  wire [1:0] n16308_o;
  wire [2:0] n16309_o;
  wire n16311_o;
  wire n16316_o;
  wire [1:0] n16317_o;
  wire n16319_o;
  wire n16320_o;
  wire n16321_o;
  wire n16322_o;
  wire n16323_o;
  wire n16324_o;
  wire n16326_o;
  wire n16328_o;
  wire n16329_o;
  wire n16330_o;
  wire [1:0] n16331_o;
  wire n16332_o;
  wire n16333_o;
  wire [1:0] n16334_o;
  reg n16335_o;
  wire [1:0] n16336_o;
  wire n16337_o;
  wire n16338_o;
  wire n16339_o;
  wire n16340_o;
  wire [16:0] n16341_o;
  wire [12:0] n16342_o;
  wire [721:0] n16343_o;
  wire n16344_o;
  wire n16345_o;
  wire n16346_o;
  wire [6:0] n16349_o;
  wire n16351_o;
  wire n16354_o;
  wire n16355_o;
  wire n16356_o;
  wire n16357_o;
  wire n16358_o;
  wire [1:0] n16359_o;
  wire n16360_o;
  wire n16361_o;
  wire n16362_o;
  wire n16363_o;
  wire n16364_o;
  wire n16365_o;
  wire n16367_o;
  wire n16368_o;
  wire n16370_o;
  wire n16371_o;
  wire n16372_o;
  wire n16373_o;
  wire n16374_o;
  wire n16375_o;
  wire n16376_o;
  wire n16378_o;
  wire n16379_o;
  wire [2:0] n16380_o;
  reg n16381_o;
  wire n16383_o;
  wire n16385_o;
  wire n16386_o;
  wire [6:0] n16387_o;
  wire n16388_o;
  wire n16389_o;
  wire n16392_o;
  wire n16394_o;
  wire n16395_o;
  wire n16396_o;
  wire n16397_o;
  wire n16398_o;
  wire n16399_o;
  wire [1:0] n16400_o;
  wire [2:0] n16402_o;
  wire n16403_o;
  wire [3:0] n16404_o;
  wire n16405_o;
  wire n16406_o;
  wire n16407_o;
  wire n16408_o;
  wire n16409_o;
  wire n16410_o;
  wire n16412_o;
  wire n16413_o;
  wire n16414_o;
  wire n16416_o;
  wire n16418_o;
  wire n16419_o;
  wire [1:0] n16422_o;
  wire n16423_o;
  wire n16424_o;
  wire n16425_o;
  wire n16426_o;
  wire n16429_o;
  wire n16431_o;
  wire [1:0] n16432_o;
  wire [2:0] n16434_o;
  wire n16435_o;
  wire [3:0] n16436_o;
  wire [79:0] n16437_o;
  wire [1:0] n16438_o;
  wire n16440_o;
  wire n16442_o;
  wire n16443_o;
  wire [2:0] n16444_o;
  wire n16447_o;
  wire n16450_o;
  wire n16451_o;
  wire n16452_o;
  wire n16454_o;
  wire n16455_o;
  wire [9:0] n16456_o;
  wire n16458_o;
  wire [12:0] n16460_o;
  wire [6:0] n16464_o;
  wire [6:0] n16465_o;
  wire [12:0] n16466_o;
  wire [6:0] n16467_o;
  wire [12:0] n16468_o;
  wire n16471_o;
  wire n16474_o;
  wire n16476_o;
  wire [12:0] n16477_o;
  wire [6:0] n16481_o;
  wire [6:0] n16482_o;
  wire [12:0] n16483_o;
  wire n16485_o;
  wire n16487_o;
  wire n16488_o;
  wire [12:0] n16491_o;
  wire [12:0] n16492_o;
  wire n16493_o;
  wire n16494_o;
  wire [6:0] n16497_o;
  wire n16500_o;
  wire [1:0] n16503_o;
  wire [6:0] n16504_o;
  wire n16505_o;
  wire n16506_o;
  wire [12:0] n16507_o;
  wire [12:0] n16508_o;
  wire n16510_o;
  wire n16513_o;
  wire n16515_o;
  wire n16517_o;
  wire n16518_o;
  wire [1:0] n16521_o;
  wire n16523_o;
  wire n16524_o;
  wire n16525_o;
  wire n16526_o;
  wire n16527_o;
  wire n16528_o;
  wire n16529_o;
  wire n16533_o;
  wire [1:0] n16534_o;
  wire [1:0] n16535_o;
  wire n16536_o;
  wire [3:0] n16538_o;
  wire [12:0] n16539_o;
  wire [12:0] n16540_o;
  wire [1:0] n16544_o;
  wire [3:0] n16546_o;
  wire [1:0] n16547_o;
  wire [14:0] n16548_o;
  wire [6:0] n16549_o;
  wire [1:0] n16550_o;
  wire [1:0] n16551_o;
  wire n16552_o;
  wire n16553_o;
  wire [1:0] n16554_o;
  wire [1:0] n16555_o;
  wire [1:0] n16556_o;
  wire [12:0] n16557_o;
  wire [12:0] n16558_o;
  wire n16561_o;
  wire n16563_o;
  wire [63:0] n16565_o;
  wire n16566_o;
  wire n16567_o;
  wire [2:0] n16568_o;
  wire n16569_o;
  wire n16577_o;
  wire [1:0] n16578_o;
  wire [2:0] n16579_o;
  wire n16580_o;
  wire [1:0] n16581_o;
  wire [2:0] n16582_o;
  wire n16583_o;
  wire [2:0] n16584_o;
  wire n16586_o;
  wire n16591_o;
  wire [1:0] n16592_o;
  wire n16594_o;
  wire n16595_o;
  wire n16596_o;
  wire n16597_o;
  wire n16598_o;
  wire n16599_o;
  wire n16601_o;
  wire n16603_o;
  wire n16604_o;
  wire n16605_o;
  wire [1:0] n16606_o;
  wire n16607_o;
  wire n16608_o;
  wire [1:0] n16609_o;
  reg n16610_o;
  wire [1:0] n16611_o;
  wire n16612_o;
  wire n16615_o;
  wire n16616_o;
  wire [6:0] n16618_o;
  wire n16621_o;
  wire n16624_o;
  wire [1:0] n16627_o;
  wire [6:0] n16628_o;
  wire [12:0] n16629_o;
  wire n16631_o;
  wire n16633_o;
  wire n16634_o;
  wire n16636_o;
  wire n16638_o;
  wire n16639_o;
  wire n16640_o;
  wire n16641_o;
  wire n16643_o;
  wire n16645_o;
  wire n16647_o;
  wire [6:0] n16649_o;
  wire n16652_o;
  wire n16653_o;
  wire n16654_o;
  wire [6:0] n16656_o;
  wire n16659_o;
  wire n16662_o;
  wire [1:0] n16665_o;
  wire [6:0] n16666_o;
  wire n16667_o;
  wire n16669_o;
  wire n16671_o;
  wire n16672_o;
  wire n16673_o;
  wire n16674_o;
  wire n16675_o;
  wire n16676_o;
  wire n16678_o;
  wire n16679_o;
  wire n16680_o;
  wire n16681_o;
  wire n16682_o;
  wire n16683_o;
  wire [12:0] n16685_o;
  wire n16687_o;
  wire [6:0] n16689_o;
  wire n16692_o;
  wire [1:0] n16695_o;
  wire [2:0] n16696_o;
  wire [6:0] n16697_o;
  wire [2:0] n16698_o;
  wire [2:0] n16699_o;
  wire [12:0] n16700_o;
  wire n16701_o;
  wire n16702_o;
  wire n16703_o;
  wire n16704_o;
  wire n16706_o;
  wire n16708_o;
  wire n16710_o;
  wire n16711_o;
  wire [79:0] n16712_o;
  wire [1:0] n16713_o;
  wire n16715_o;
  wire n16716_o;
  wire n16717_o;
  wire n16718_o;
  wire n16719_o;
  wire n16720_o;
  wire [79:0] n16721_o;
  wire [1:0] n16722_o;
  wire n16724_o;
  wire n16725_o;
  wire n16726_o;
  wire n16727_o;
  wire n16728_o;
  wire n16729_o;
  wire n16730_o;
  wire [79:0] n16731_o;
  wire [1:0] n16732_o;
  wire n16734_o;
  wire n16735_o;
  wire n16736_o;
  wire n16737_o;
  wire n16738_o;
  wire n16739_o;
  wire n16741_o;
  wire n16742_o;
  wire n16745_o;
  wire n16746_o;
  wire [79:0] n16747_o;
  wire [1:0] n16748_o;
  wire n16750_o;
  wire n16751_o;
  wire n16753_o;
  wire [79:0] n16754_o;
  wire [1:0] n16755_o;
  wire n16757_o;
  wire n16758_o;
  wire n16760_o;
  wire [79:0] n16761_o;
  wire [1:0] n16762_o;
  wire n16764_o;
  wire n16765_o;
  wire [1:0] n16767_o;
  wire [1:0] n16768_o;
  wire [1:0] n16769_o;
  wire n16772_o;
  wire [1:0] n16773_o;
  wire [79:0] n16774_o;
  wire n16775_o;
  wire n16776_o;
  wire n16777_o;
  wire [79:0] n16778_o;
  wire [12:0] n16779_o;
  wire [79:0] n16780_o;
  wire [1:0] n16781_o;
  wire n16783_o;
  wire [79:0] n16784_o;
  wire n16785_o;
  wire n16786_o;
  wire n16787_o;
  wire [79:0] n16788_o;
  wire [12:0] n16789_o;
  wire [79:0] n16790_o;
  wire [1:0] n16791_o;
  wire n16793_o;
  wire [79:0] n16794_o;
  wire n16795_o;
  wire n16796_o;
  wire n16797_o;
  wire [79:0] n16798_o;
  wire [12:0] n16799_o;
  wire [79:0] n16800_o;
  wire [1:0] n16801_o;
  wire [1:0] n16802_o;
  reg n16803_o;
  reg [1:0] n16804_o;
  reg [12:0] n16805_o;
  wire n16807_o;
  wire [79:0] n16808_o;
  reg [1:0] n16814_o;
  reg [1:0] n16836_o;
  reg [1:0] n16843_o;
  reg n16847_o;
  reg n16852_o;
  reg n16857_o;
  reg n16862_o;
  wire n16864_o;
  wire n16868_o;
  wire n16869_o;
  reg n16872_o;
  wire [2:0] n16873_o;
  wire [2:0] n16877_o;
  wire [2:0] n16878_o;
  reg [2:0] n16881_o;
  reg n16885_o;
  reg [1:0] n16899_o;
  reg [1:0] n16915_o;
  reg [1:0] n16925_o;
  reg n16934_o;
  reg [6:0] n16937_o;
  reg n16939_o;
  wire n16940_o;
  wire n16941_o;
  wire n16942_o;
  wire n16943_o;
  wire n16944_o;
  reg n16946_o;
  wire n16947_o;
  wire n16948_o;
  wire n16949_o;
  wire n16950_o;
  wire n16951_o;
  reg n16953_o;
  wire n16954_o;
  wire n16955_o;
  wire n16956_o;
  wire n16957_o;
  reg n16959_o;
  wire n16960_o;
  wire n16961_o;
  wire n16962_o;
  wire n16963_o;
  wire n16964_o;
  reg n16966_o;
  wire n16967_o;
  wire n16968_o;
  wire n16969_o;
  wire n16970_o;
  wire n16971_o;
  reg n16973_o;
  wire n16974_o;
  wire n16975_o;
  wire n16976_o;
  wire n16977_o;
  wire n16978_o;
  reg n16980_o;
  wire n16981_o;
  wire n16982_o;
  wire n16983_o;
  wire n16984_o;
  wire n16985_o;
  reg n16987_o;
  wire n16988_o;
  wire n16989_o;
  wire n16990_o;
  wire n16991_o;
  wire n16992_o;
  reg n16994_o;
  wire n16995_o;
  wire n16996_o;
  wire n16997_o;
  wire n16998_o;
  reg n17000_o;
  wire n17001_o;
  wire n17002_o;
  wire n17003_o;
  wire n17004_o;
  reg n17006_o;
  wire n17007_o;
  wire n17008_o;
  wire n17009_o;
  wire n17010_o;
  reg n17012_o;
  wire n17013_o;
  wire n17014_o;
  wire n17015_o;
  wire n17016_o;
  reg n17018_o;
  wire n17019_o;
  wire n17020_o;
  wire n17021_o;
  wire n17022_o;
  wire n17023_o;
  wire n17024_o;
  reg n17026_o;
  wire n17027_o;
  wire n17028_o;
  wire n17029_o;
  wire n17030_o;
  wire n17031_o;
  wire n17032_o;
  reg n17034_o;
  wire n17035_o;
  wire n17036_o;
  wire n17037_o;
  wire n17038_o;
  wire n17039_o;
  wire n17040_o;
  reg n17042_o;
  wire n17043_o;
  wire n17044_o;
  wire n17045_o;
  wire n17046_o;
  wire n17047_o;
  wire n17048_o;
  reg n17050_o;
  wire n17051_o;
  wire n17052_o;
  wire n17053_o;
  wire n17054_o;
  reg n17056_o;
  wire n17057_o;
  wire n17058_o;
  wire n17059_o;
  wire n17060_o;
  wire n17061_o;
  wire n17062_o;
  wire n17063_o;
  reg n17065_o;
  wire n17066_o;
  wire n17067_o;
  wire n17068_o;
  wire n17069_o;
  wire n17070_o;
  wire n17071_o;
  wire n17072_o;
  reg n17074_o;
  wire n17075_o;
  wire n17076_o;
  wire n17077_o;
  wire n17078_o;
  reg n17080_o;
  wire n17081_o;
  wire n17082_o;
  wire n17083_o;
  wire n17084_o;
  reg n17086_o;
  wire n17087_o;
  wire n17088_o;
  wire n17089_o;
  wire n17090_o;
  wire n17091_o;
  reg n17093_o;
  wire n17094_o;
  wire n17095_o;
  wire n17096_o;
  wire n17097_o;
  wire n17098_o;
  reg n17100_o;
  wire n17101_o;
  wire n17102_o;
  wire n17103_o;
  wire n17104_o;
  reg n17106_o;
  wire n17107_o;
  wire n17108_o;
  wire n17109_o;
  wire n17110_o;
  reg n17112_o;
  wire n17113_o;
  wire n17114_o;
  wire n17115_o;
  wire n17116_o;
  reg n17118_o;
  wire n17119_o;
  wire n17120_o;
  wire n17121_o;
  wire n17122_o;
  reg n17124_o;
  wire n17125_o;
  wire n17126_o;
  wire n17127_o;
  wire n17128_o;
  reg n17130_o;
  wire n17131_o;
  wire n17132_o;
  wire n17133_o;
  wire n17134_o;
  reg n17136_o;
  wire n17137_o;
  wire n17138_o;
  wire n17139_o;
  wire n17140_o;
  reg n17142_o;
  wire n17143_o;
  wire n17144_o;
  wire n17145_o;
  wire n17146_o;
  reg n17148_o;
  wire n17149_o;
  wire n17150_o;
  wire n17151_o;
  wire n17152_o;
  reg n17154_o;
  wire n17155_o;
  reg n17157_o;
  wire n17158_o;
  wire n17159_o;
  wire n17160_o;
  reg n17162_o;
  wire [1:0] n17163_o;
  wire [1:0] n17164_o;
  wire [1:0] n17165_o;
  reg [1:0] n17167_o;
  wire [12:0] n17168_o;
  wire [12:0] n17169_o;
  reg [12:0] n17171_o;
  wire [12:0] n17172_o;
  reg [12:0] n17174_o;
  reg n17176_o;
  reg n17178_o;
  wire n17179_o;
  wire n17180_o;
  wire n17181_o;
  wire n17182_o;
  reg n17184_o;
  wire n17185_o;
  wire n17186_o;
  wire n17187_o;
  wire n17188_o;
  reg n17190_o;
  wire n17191_o;
  wire n17192_o;
  wire n17193_o;
  wire n17194_o;
  reg n17196_o;
  wire n17197_o;
  wire n17198_o;
  wire n17199_o;
  wire n17200_o;
  reg n17202_o;
  reg [4:0] n17204_o;
  wire n17205_o;
  wire n17206_o;
  wire n17207_o;
  reg n17209_o;
  wire n17210_o;
  wire n17211_o;
  wire n17212_o;
  reg n17214_o;
  wire n17215_o;
  wire n17216_o;
  wire n17217_o;
  reg n17219_o;
  wire [2:0] n17220_o;
  wire [2:0] n17221_o;
  wire [2:0] n17222_o;
  reg [2:0] n17224_o;
  wire n17225_o;
  wire n17226_o;
  wire n17227_o;
  reg n17229_o;
  wire n17230_o;
  wire n17231_o;
  wire n17232_o;
  reg n17234_o;
  wire n17235_o;
  wire n17236_o;
  wire n17237_o;
  reg n17239_o;
  wire n17240_o;
  wire n17241_o;
  wire n17242_o;
  wire n17243_o;
  reg n17245_o;
  wire n17246_o;
  wire n17247_o;
  wire n17248_o;
  wire n17249_o;
  reg n17251_o;
  wire n17252_o;
  wire n17253_o;
  reg n17255_o;
  wire [1:0] n17256_o;
  wire [1:0] n17257_o;
  reg [1:0] n17259_o;
  reg [1:0] n17261_o;
  reg [1:0] n17263_o;
  wire n17264_o;
  reg n17266_o;
  wire n17267_o;
  reg n17269_o;
  wire n17270_o;
  reg n17272_o;
  wire n17273_o;
  reg n17275_o;
  wire n17276_o;
  reg n17278_o;
  reg n17280_o;
  wire [119:0] n17313_o;
  wire [127:0] n17315_o;
  wire n17338_o;
  wire n17339_o;
  wire n17340_o;
  wire [3:0] n17351_o;
  reg [3:0] n17354_o;
  wire [3:0] n17355_o;
  reg [3:0] n17358_o;
  wire [3:0] n17359_o;
  reg [3:0] n17362_o;
  wire [3:0] n17363_o;
  reg [3:0] n17366_o;
  wire [3:0] n17367_o;
  reg [3:0] n17370_o;
  wire [3:0] n17371_o;
  reg [3:0] n17374_o;
  wire [3:0] n17375_o;
  reg [3:0] n17378_o;
  wire [3:0] n17379_o;
  reg [3:0] n17382_o;
  reg n17393_o;
  reg n17407_o;
  reg n17415_o;
  reg n17420_o;
  reg n17424_o;
  reg n17433_o;
  reg n17442_o;
  reg n17454_o;
  reg n17459_o;
  reg n17464_o;
  reg n17468_o;
  reg n17476_o;
  reg n17480_o;
  reg n17493_o;
  reg n17497_o;
  reg n17504_o;
  wire n17509_o;
  wire [1:0] n17513_o;
  wire [3:0] n17515_o;
  wire [3:0] n17516_o;
  wire [2:0] n17517_o;
  wire [2:0] n17518_o;
  wire [2:0] n17519_o;
  wire n17521_o;
  wire n17523_o;
  wire n17525_o;
  wire [721:0] n17526_o;
  wire n17527_o;
  wire n17528_o;
  wire n17529_o;
  wire n17530_o;
  wire n17531_o;
  wire n17532_o;
  wire n17533_o;
  wire n17534_o;
  wire n17537_o;
  wire n17538_o;
  wire [6:0] n17541_o;
  wire n17542_o;
  wire n17543_o;
  wire n17544_o;
  wire n17546_o;
  wire [61:0] n17547_o;
  wire [63:0] n17549_o;
  wire n17551_o;
  wire [61:0] n17552_o;
  wire [63:0] n17554_o;
  wire n17556_o;
  wire [63:0] n17557_o;
  wire n17559_o;
  wire [61:0] n17560_o;
  wire [63:0] n17562_o;
  wire [2:0] n17563_o;
  reg [63:0] n17564_o;
  wire [61:0] n17565_o;
  wire [63:0] n17567_o;
  wire n17569_o;
  wire [26:0] n17571_o;
  wire [27:0] n17573_o;
  wire [63:0] n17575_o;
  wire n17577_o;
  wire [63:0] n17578_o;
  wire n17580_o;
  wire [61:0] n17581_o;
  wire [63:0] n17583_o;
  wire [2:0] n17584_o;
  reg [63:0] n17585_o;
  wire n17586_o;
  wire n17587_o;
  wire [1:0] n17591_o;
  wire n17593_o;
  wire n17595_o;
  wire [79:0] n17596_o;
  wire [63:0] n17597_o;
  wire n17599_o;
  wire [63:0] n17600_o;
  wire [69:0] n17602_o;
  wire [55:0] n17603_o;
  wire [125:0] n17604_o;
  wire [127:0] n17606_o;
  wire n17608_o;
  wire [2:0] n17609_o;
  wire [57:0] n17610_o;
  reg [57:0] n17612_o;
  wire [52:0] n17613_o;
  wire [52:0] n17614_o;
  reg [52:0] n17616_o;
  wire [1:0] n17617_o;
  wire [1:0] n17618_o;
  reg [1:0] n17620_o;
  wire n17621_o;
  wire n17622_o;
  reg n17624_o;
  wire [7:0] n17625_o;
  wire [7:0] n17626_o;
  reg [7:0] n17628_o;
  wire [5:0] n17629_o;
  reg [5:0] n17631_o;
  wire [127:0] n17638_o;
  wire [127:0] n17639_o;
  wire [127:0] n17640_o;
  wire [127:0] n17641_o;
  wire [63:0] n17642_o;
  wire [63:0] n17643_o;
  wire [63:0] n17644_o;
  wire [63:0] n17645_o;
  wire n17646_o;
  wire n17647_o;
  wire [63:0] n17648_o;
  wire [63:0] n17649_o;
  wire [63:0] n17650_o;
  wire [63:0] n17651_o;
  wire n17652_o;
  wire [12:0] n17653_o;
  wire [12:0] n17655_o;
  wire [12:0] n17656_o;
  wire [12:0] n17657_o;
  wire n17659_o;
  wire n17661_o;
  wire [5:0] n17663_o;
  wire n17670_o;
  wire n17673_o;
  localparam [63:0] n17674_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire n17677_o;
  wire n17679_o;
  wire n17680_o;
  wire n17683_o;
  wire n17685_o;
  wire n17686_o;
  wire n17689_o;
  wire n17691_o;
  wire n17692_o;
  wire n17695_o;
  wire n17697_o;
  wire n17698_o;
  wire n17701_o;
  wire n17703_o;
  wire n17704_o;
  wire n17707_o;
  wire n17709_o;
  wire n17710_o;
  wire n17713_o;
  wire n17715_o;
  wire n17716_o;
  wire n17719_o;
  wire n17721_o;
  wire n17722_o;
  wire n17725_o;
  wire n17727_o;
  wire n17728_o;
  wire n17731_o;
  wire n17733_o;
  wire n17734_o;
  wire n17737_o;
  wire n17739_o;
  wire n17740_o;
  wire n17743_o;
  wire n17745_o;
  wire n17746_o;
  wire n17749_o;
  wire n17751_o;
  wire n17752_o;
  wire n17755_o;
  wire n17757_o;
  wire n17758_o;
  wire n17761_o;
  wire n17763_o;
  wire n17764_o;
  wire n17767_o;
  wire n17769_o;
  wire n17770_o;
  wire n17773_o;
  wire n17775_o;
  wire n17776_o;
  wire n17779_o;
  wire n17781_o;
  wire n17782_o;
  wire n17785_o;
  wire n17787_o;
  wire n17788_o;
  wire n17791_o;
  wire n17793_o;
  wire n17794_o;
  wire n17797_o;
  wire n17799_o;
  wire n17800_o;
  wire n17803_o;
  wire n17805_o;
  wire n17806_o;
  wire n17809_o;
  wire n17811_o;
  wire n17812_o;
  wire n17815_o;
  wire n17817_o;
  wire n17818_o;
  wire n17821_o;
  wire n17823_o;
  wire n17824_o;
  wire n17827_o;
  wire n17829_o;
  wire n17830_o;
  wire n17833_o;
  wire n17835_o;
  wire n17836_o;
  wire n17839_o;
  wire n17841_o;
  wire n17842_o;
  wire n17845_o;
  wire n17847_o;
  wire n17848_o;
  wire n17851_o;
  wire n17853_o;
  wire n17854_o;
  wire n17857_o;
  wire n17859_o;
  wire n17860_o;
  wire n17863_o;
  wire n17865_o;
  wire n17866_o;
  wire n17869_o;
  wire n17871_o;
  wire n17872_o;
  wire n17875_o;
  wire n17877_o;
  wire n17878_o;
  wire n17881_o;
  wire n17883_o;
  wire n17884_o;
  wire n17887_o;
  wire n17889_o;
  wire n17890_o;
  wire n17893_o;
  wire n17895_o;
  wire n17896_o;
  wire n17899_o;
  wire n17901_o;
  wire n17902_o;
  wire n17905_o;
  wire n17907_o;
  wire n17908_o;
  wire n17911_o;
  wire n17913_o;
  wire n17914_o;
  wire n17917_o;
  wire n17919_o;
  wire n17920_o;
  wire n17923_o;
  wire n17925_o;
  wire n17926_o;
  wire n17929_o;
  wire n17931_o;
  wire n17932_o;
  wire n17935_o;
  wire n17937_o;
  wire n17938_o;
  wire n17941_o;
  wire n17943_o;
  wire n17944_o;
  wire n17947_o;
  wire n17949_o;
  wire n17950_o;
  wire n17953_o;
  wire n17955_o;
  wire n17956_o;
  wire n17959_o;
  wire n17961_o;
  wire n17962_o;
  wire n17965_o;
  wire n17967_o;
  wire n17968_o;
  wire n17971_o;
  wire n17973_o;
  wire n17974_o;
  wire n17977_o;
  wire n17979_o;
  wire n17980_o;
  wire n17983_o;
  wire n17985_o;
  wire n17986_o;
  wire n17989_o;
  wire n17991_o;
  wire n17992_o;
  wire n17995_o;
  wire n17997_o;
  wire n17998_o;
  wire n18001_o;
  wire n18003_o;
  wire n18004_o;
  wire n18007_o;
  wire n18009_o;
  wire n18010_o;
  wire n18013_o;
  wire n18015_o;
  wire n18016_o;
  wire n18019_o;
  wire n18021_o;
  wire n18022_o;
  wire n18025_o;
  wire n18027_o;
  wire n18028_o;
  wire n18031_o;
  wire n18033_o;
  wire n18034_o;
  wire n18037_o;
  wire n18039_o;
  wire n18040_o;
  wire n18043_o;
  wire n18045_o;
  wire n18046_o;
  wire n18047_o;
  wire n18049_o;
  wire n18051_o;
  wire [63:0] n18052_o;
  wire [63:0] n18054_o;
  wire [63:0] n18056_o;
  wire [1:0] n18057_o;
  wire [63:0] n18058_o;
  wire n18060_o;
  wire [79:0] n18061_o;
  wire [63:0] n18062_o;
  wire n18064_o;
  wire [79:0] n18065_o;
  wire [63:0] n18066_o;
  wire n18068_o;
  wire [79:0] n18069_o;
  wire [63:0] n18070_o;
  wire [2:0] n18071_o;
  reg [63:0] n18072_o;
  wire [63:0] n18073_o;
  wire n18074_o;
  wire n18075_o;
  wire n18077_o;
  wire [63:0] n18078_o;
  wire [63:0] n18079_o;
  wire n18081_o;
  wire [63:0] n18082_o;
  wire n18084_o;
  wire n18085_o;
  wire n18086_o;
  wire n18087_o;
  wire [3:0] n18150_o;
  wire [3:0] n18151_o;
  wire [3:0] n18152_o;
  wire [3:0] n18153_o;
  wire [3:0] n18154_o;
  wire [3:0] n18155_o;
  wire [3:0] n18156_o;
  wire [3:0] n18157_o;
  wire [3:0] n18158_o;
  wire [3:0] n18159_o;
  wire [3:0] n18160_o;
  wire [3:0] n18161_o;
  wire [3:0] n18162_o;
  wire [3:0] n18163_o;
  wire [3:0] n18164_o;
  wire [3:0] n18165_o;
  wire [15:0] n18166_o;
  wire [15:0] n18167_o;
  wire [15:0] n18168_o;
  wire [15:0] n18169_o;
  wire [63:0] n18170_o;
  wire n18172_o;
  wire [5:0] n18173_o;
  wire [63:0] n18174_o;
  wire [2:0] n18175_o;
  reg [63:0] n18177_o;
  wire [63:0] n18179_o;
  wire [63:0] n18180_o;
  wire [12:0] n18181_o;
  wire n18183_o;
  wire [12:0] n18184_o;
  wire n18186_o;
  wire n18187_o;
  wire [63:0] n18189_o;
  wire n18190_o;
  wire n18191_o;
  wire [64:0] n18192_o;
  wire [54:0] n18193_o;
  wire [119:0] n18194_o;
  wire [6:0] n18195_o;
  wire [1:0] n18203_o;
  wire [94:0] n18204_o;
  wire n18206_o;
  wire [87:0] n18207_o;
  wire [94:0] n18209_o;
  wire n18211_o;
  wire [30:0] n18212_o;
  wire [94:0] n18214_o;
  wire n18216_o;
  wire [62:0] n18217_o;
  wire [94:0] n18219_o;
  wire [2:0] n18220_o;
  reg [94:0] n18221_o;
  wire [1:0] n18223_o;
  wire [70:0] n18224_o;
  wire n18226_o;
  wire [70:0] n18227_o;
  wire n18229_o;
  wire [70:0] n18230_o;
  wire n18232_o;
  wire [70:0] n18233_o;
  wire [2:0] n18234_o;
  reg [70:0] n18235_o;
  wire [2:0] n18237_o;
  wire [63:0] n18238_o;
  wire n18240_o;
  wire [63:0] n18241_o;
  wire n18243_o;
  wire [63:0] n18244_o;
  wire n18246_o;
  wire [63:0] n18247_o;
  wire n18249_o;
  wire [63:0] n18250_o;
  wire n18252_o;
  wire [63:0] n18253_o;
  wire n18255_o;
  wire [63:0] n18256_o;
  wire n18258_o;
  wire [63:0] n18259_o;
  wire [6:0] n18260_o;
  reg [63:0] n18261_o;
  wire [63:0] n18264_o;
  wire [63:0] n18265_o;
  wire [63:0] n18266_o;
  wire [63:0] n18267_o;
  wire n18269_o;
  wire [28:0] n18271_o;
  wire [28:0] n18272_o;
  wire [30:0] n18273_o;
  wire [30:0] n18274_o;
  wire [30:0] n18275_o;
  wire [32:0] n18276_o;
  wire [63:0] n18277_o;
  wire n18279_o;
  wire n18281_o;
  wire [63:0] n18282_o;
  wire n18284_o;
  wire [31:0] n18285_o;
  wire [31:0] n18286_o;
  wire [31:0] n18287_o;
  wire [63:0] n18289_o;
  wire n18291_o;
  wire n18293_o;
  wire n18295_o;
  wire n18297_o;
  wire [31:0] n18298_o;
  wire [31:0] n18299_o;
  wire [63:0] n18300_o;
  wire n18302_o;
  wire [31:0] n18303_o;
  wire [31:0] n18304_o;
  wire [63:0] n18305_o;
  wire n18307_o;
  wire [28:0] n18309_o;
  wire [63:0] n18311_o;
  wire n18313_o;
  wire n18315_o;
  wire n18317_o;
  wire n18319_o;
  wire n18321_o;
  wire n18323_o;
  wire n18325_o;
  wire n18327_o;
  wire n18329_o;
  wire [14:0] n18330_o;
  reg [63:0] n18343_o;
  wire [2:0] n18344_o;
  reg [63:0] n18345_o;
  wire [55:0] n18347_o;
  wire [55:0] n18348_o;
  wire [55:0] n18349_o;
  wire n18350_o;
  wire n18351_o;
  wire [55:0] n18352_o;
  wire [55:0] n18353_o;
  wire n18355_o;
  wire [55:0] n18356_o;
  wire n18358_o;
  wire [55:0] n18359_o;
  wire [7:0] n18360_o;
  wire n18362_o;
  wire n18364_o;
  wire n18366_o;
  wire [2:0] n18368_o;
  reg [55:0] n18369_o;
  reg n18370_o;
  wire [56:0] n18371_o;
  wire [56:0] n18372_o;
  wire [56:0] n18373_o;
  wire [76:0] n18374_o;
  wire [76:0] n18375_o;
  wire [76:0] n18376_o;
  wire [76:0] n18377_o;
  wire [76:0] n18378_o;
  wire [2:0] n18382_o;
  wire [2:0] n18383_o;
  wire [2:0] n18384_o;
  wire [76:0] n18385_o;
  wire [76:0] n18386_o;
  wire [76:0] n18387_o;
  wire [76:0] n18388_o;
  wire [76:0] n18389_o;
  wire [2:0] n18393_o;
  wire [2:0] n18394_o;
  wire [2:0] n18395_o;
  wire [76:0] n18396_o;
  wire [76:0] n18397_o;
  wire [76:0] n18398_o;
  wire [76:0] n18399_o;
  wire [76:0] n18400_o;
  wire [2:0] n18401_o;
  wire [2:0] n18402_o;
  wire [2:0] n18403_o;
  wire n18405_o;
  wire [12:0] n18406_o;
  wire [63:0] n18408_o;
  wire n18420_o;
  wire n18423_o;
  wire n18425_o;
  wire n18427_o;
  wire n18429_o;
  wire n18431_o;
  wire n18433_o;
  wire n18435_o;
  wire n18437_o;
  wire n18439_o;
  wire n18441_o;
  wire n18443_o;
  wire n18445_o;
  wire n18447_o;
  wire n18449_o;
  wire n18451_o;
  wire n18453_o;
  wire n18455_o;
  wire n18457_o;
  wire n18459_o;
  wire n18461_o;
  wire n18463_o;
  wire n18465_o;
  wire n18467_o;
  wire n18469_o;
  wire n18471_o;
  wire n18473_o;
  wire n18475_o;
  wire n18477_o;
  wire n18479_o;
  wire n18481_o;
  wire n18483_o;
  wire n18485_o;
  wire n18487_o;
  wire n18489_o;
  wire n18491_o;
  wire n18493_o;
  wire n18495_o;
  wire n18497_o;
  wire n18499_o;
  wire n18501_o;
  wire n18503_o;
  wire n18505_o;
  wire n18507_o;
  wire n18509_o;
  wire n18511_o;
  wire n18513_o;
  wire n18515_o;
  wire n18517_o;
  wire n18519_o;
  wire n18521_o;
  wire n18523_o;
  wire n18525_o;
  wire n18527_o;
  wire n18529_o;
  wire n18531_o;
  wire n18533_o;
  wire n18535_o;
  wire n18537_o;
  wire n18539_o;
  wire n18541_o;
  wire n18543_o;
  wire n18545_o;
  wire n18547_o;
  wire [63:0] n18548_o;
  wire [63:0] n18561_o;
  wire [63:0] n18563_o;
  wire [63:0] n18565_o;
  wire n18576_o;
  wire n18577_o;
  wire n18578_o;
  wire n18579_o;
  wire n18581_o;
  wire n18583_o;
  wire n18584_o;
  wire n18585_o;
  wire n18586_o;
  wire n18587_o;
  wire n18588_o;
  wire n18589_o;
  wire n18590_o;
  wire n18591_o;
  wire n18592_o;
  wire n18593_o;
  wire n18594_o;
  wire n18595_o;
  wire n18596_o;
  wire n18597_o;
  wire n18598_o;
  wire n18599_o;
  wire n18600_o;
  wire n18601_o;
  wire n18602_o;
  wire n18603_o;
  wire n18604_o;
  wire n18605_o;
  wire n18606_o;
  wire n18607_o;
  wire n18608_o;
  wire n18609_o;
  wire n18610_o;
  wire n18611_o;
  wire n18612_o;
  wire n18613_o;
  wire n18614_o;
  wire n18615_o;
  wire n18616_o;
  wire n18617_o;
  wire n18618_o;
  wire n18619_o;
  wire n18620_o;
  wire n18621_o;
  wire n18622_o;
  wire n18623_o;
  wire n18624_o;
  wire n18625_o;
  wire n18626_o;
  wire n18627_o;
  wire n18628_o;
  wire n18629_o;
  wire n18630_o;
  wire n18631_o;
  wire n18632_o;
  wire n18633_o;
  wire n18634_o;
  wire n18635_o;
  wire n18636_o;
  wire n18637_o;
  wire n18638_o;
  wire n18639_o;
  wire n18640_o;
  wire n18641_o;
  wire n18642_o;
  wire n18643_o;
  wire n18644_o;
  wire n18645_o;
  wire n18646_o;
  wire n18647_o;
  wire n18648_o;
  wire n18649_o;
  wire n18650_o;
  wire n18651_o;
  wire n18652_o;
  wire n18653_o;
  wire n18654_o;
  wire n18655_o;
  wire n18656_o;
  wire n18657_o;
  wire n18658_o;
  wire n18659_o;
  wire n18660_o;
  wire n18661_o;
  wire n18662_o;
  wire n18663_o;
  wire n18664_o;
  wire n18665_o;
  wire n18666_o;
  wire n18667_o;
  wire n18668_o;
  wire n18669_o;
  wire n18670_o;
  wire n18671_o;
  wire n18672_o;
  wire n18673_o;
  wire n18674_o;
  wire n18675_o;
  wire n18676_o;
  wire n18677_o;
  wire n18678_o;
  wire n18679_o;
  wire n18680_o;
  wire n18681_o;
  wire n18682_o;
  wire n18683_o;
  wire n18684_o;
  wire n18685_o;
  wire n18686_o;
  wire n18687_o;
  wire n18688_o;
  wire n18689_o;
  wire n18690_o;
  wire n18691_o;
  wire n18692_o;
  wire n18693_o;
  wire n18694_o;
  wire n18695_o;
  wire n18696_o;
  wire n18697_o;
  wire n18698_o;
  wire n18699_o;
  wire n18700_o;
  wire n18701_o;
  wire n18702_o;
  wire n18703_o;
  wire n18704_o;
  wire n18705_o;
  wire n18706_o;
  wire n18707_o;
  wire n18708_o;
  wire n18709_o;
  wire n18710_o;
  wire n18711_o;
  wire n18712_o;
  wire n18713_o;
  wire n18714_o;
  wire n18715_o;
  wire n18716_o;
  wire n18717_o;
  wire n18718_o;
  wire n18719_o;
  wire n18720_o;
  wire n18721_o;
  wire n18722_o;
  wire n18723_o;
  wire n18724_o;
  wire n18725_o;
  wire n18726_o;
  wire n18727_o;
  wire n18728_o;
  wire n18729_o;
  wire n18730_o;
  wire n18731_o;
  wire n18732_o;
  wire n18733_o;
  wire n18734_o;
  wire n18735_o;
  wire n18736_o;
  wire n18737_o;
  wire n18740_o;
  wire n18741_o;
  wire n18742_o;
  wire n18743_o;
  wire n18745_o;
  wire n18747_o;
  wire n18748_o;
  wire n18749_o;
  wire n18750_o;
  wire n18751_o;
  wire n18752_o;
  wire n18753_o;
  wire n18754_o;
  wire n18755_o;
  wire n18756_o;
  wire n18757_o;
  wire n18758_o;
  wire n18759_o;
  wire n18760_o;
  wire n18761_o;
  wire n18762_o;
  wire n18763_o;
  wire n18764_o;
  wire n18765_o;
  wire n18766_o;
  wire n18767_o;
  wire n18768_o;
  wire n18769_o;
  wire n18770_o;
  wire n18771_o;
  wire n18772_o;
  wire n18773_o;
  wire n18774_o;
  wire n18775_o;
  wire n18776_o;
  wire n18777_o;
  wire n18778_o;
  wire n18779_o;
  wire n18780_o;
  wire n18781_o;
  wire n18782_o;
  wire n18783_o;
  wire n18784_o;
  wire n18785_o;
  wire n18786_o;
  wire n18787_o;
  wire n18788_o;
  wire n18789_o;
  wire n18790_o;
  wire n18791_o;
  wire n18792_o;
  wire n18793_o;
  wire n18794_o;
  wire n18795_o;
  wire n18796_o;
  wire n18797_o;
  wire n18798_o;
  wire n18799_o;
  wire n18800_o;
  wire n18801_o;
  wire n18802_o;
  wire n18803_o;
  wire n18804_o;
  wire n18805_o;
  wire n18806_o;
  wire n18807_o;
  wire n18808_o;
  wire n18809_o;
  wire n18810_o;
  wire n18811_o;
  wire n18812_o;
  wire n18813_o;
  wire n18814_o;
  wire n18815_o;
  wire n18816_o;
  wire n18817_o;
  wire n18818_o;
  wire n18819_o;
  wire n18820_o;
  wire n18821_o;
  wire n18823_o;
  wire n18824_o;
  wire n18825_o;
  wire n18826_o;
  wire n18828_o;
  wire n18830_o;
  wire n18831_o;
  wire n18832_o;
  wire n18833_o;
  wire n18834_o;
  wire n18835_o;
  wire n18836_o;
  wire n18837_o;
  wire n18838_o;
  wire n18839_o;
  wire n18840_o;
  wire n18841_o;
  wire n18842_o;
  wire n18843_o;
  wire n18844_o;
  wire n18845_o;
  wire n18846_o;
  wire n18847_o;
  wire n18848_o;
  wire n18849_o;
  wire n18850_o;
  wire n18851_o;
  wire n18852_o;
  wire n18853_o;
  wire n18854_o;
  wire n18855_o;
  wire n18856_o;
  wire n18857_o;
  wire n18858_o;
  wire n18859_o;
  wire n18860_o;
  wire n18861_o;
  wire n18862_o;
  wire n18863_o;
  wire n18864_o;
  wire n18866_o;
  wire n18867_o;
  wire n18868_o;
  wire n18869_o;
  wire n18871_o;
  wire n18873_o;
  wire n18874_o;
  wire n18875_o;
  wire n18876_o;
  wire n18877_o;
  wire n18878_o;
  wire n18879_o;
  wire n18880_o;
  wire n18881_o;
  wire n18882_o;
  wire n18883_o;
  wire n18884_o;
  wire n18885_o;
  wire n18886_o;
  wire n18887_o;
  wire n18889_o;
  wire n18890_o;
  wire n18891_o;
  wire n18892_o;
  wire n18894_o;
  wire n18896_o;
  wire n18897_o;
  wire n18898_o;
  wire n18899_o;
  wire n18900_o;
  wire n18902_o;
  wire n18903_o;
  wire n18904_o;
  wire n18905_o;
  wire n18907_o;
  wire [5:0] n18909_o;
  wire n18920_o;
  wire n18921_o;
  wire n18923_o;
  wire n18925_o;
  wire n18926_o;
  wire n18927_o;
  wire n18928_o;
  wire n18929_o;
  wire n18930_o;
  wire n18931_o;
  wire n18932_o;
  wire n18933_o;
  wire n18934_o;
  wire n18935_o;
  wire n18936_o;
  wire n18937_o;
  wire n18938_o;
  wire n18939_o;
  wire n18940_o;
  wire n18941_o;
  wire n18942_o;
  wire n18943_o;
  wire n18944_o;
  wire n18945_o;
  wire n18946_o;
  wire n18947_o;
  wire n18948_o;
  wire n18949_o;
  wire n18950_o;
  wire n18951_o;
  wire n18952_o;
  wire n18953_o;
  wire n18954_o;
  wire n18955_o;
  wire n18956_o;
  wire n18957_o;
  wire n18958_o;
  wire n18959_o;
  wire n18960_o;
  wire n18961_o;
  wire n18962_o;
  wire n18963_o;
  wire n18964_o;
  wire n18965_o;
  wire n18966_o;
  wire n18967_o;
  wire n18968_o;
  wire n18969_o;
  wire n18970_o;
  wire n18971_o;
  wire n18972_o;
  wire n18973_o;
  wire n18974_o;
  wire n18975_o;
  wire n18976_o;
  wire n18977_o;
  wire n18978_o;
  wire n18979_o;
  wire n18980_o;
  wire n18981_o;
  wire n18982_o;
  wire n18983_o;
  wire n18984_o;
  wire n18985_o;
  wire n18986_o;
  wire n18987_o;
  wire n18988_o;
  wire n18989_o;
  wire n18990_o;
  wire n18991_o;
  wire n18992_o;
  wire n18993_o;
  wire n18994_o;
  wire n18995_o;
  wire n18996_o;
  wire n18997_o;
  wire n18998_o;
  wire n18999_o;
  wire n19000_o;
  wire n19001_o;
  wire n19002_o;
  wire n19003_o;
  wire n19004_o;
  wire n19005_o;
  wire n19006_o;
  wire n19007_o;
  wire n19008_o;
  wire n19009_o;
  wire n19010_o;
  wire n19011_o;
  wire n19012_o;
  wire n19013_o;
  wire n19014_o;
  wire n19015_o;
  wire n19016_o;
  wire n19017_o;
  wire [1:0] n19020_o;
  wire n19021_o;
  wire n19023_o;
  wire [1:0] n19025_o;
  wire n19026_o;
  wire n19027_o;
  wire [1:0] n19028_o;
  wire n19029_o;
  wire n19030_o;
  wire [1:0] n19031_o;
  wire n19032_o;
  wire n19033_o;
  wire [1:0] n19034_o;
  wire n19035_o;
  wire n19036_o;
  wire [1:0] n19037_o;
  wire n19038_o;
  wire n19039_o;
  wire [1:0] n19040_o;
  wire n19041_o;
  wire n19042_o;
  wire [1:0] n19043_o;
  wire n19044_o;
  wire n19045_o;
  wire [1:0] n19046_o;
  wire n19047_o;
  wire n19048_o;
  wire [1:0] n19049_o;
  wire n19050_o;
  wire n19051_o;
  wire [1:0] n19052_o;
  wire n19053_o;
  wire n19054_o;
  wire [1:0] n19055_o;
  wire n19056_o;
  wire n19057_o;
  wire [1:0] n19058_o;
  wire n19059_o;
  wire n19060_o;
  wire [1:0] n19061_o;
  wire n19062_o;
  wire n19063_o;
  wire [1:0] n19064_o;
  wire n19065_o;
  wire n19066_o;
  wire [1:0] n19067_o;
  wire n19068_o;
  wire n19069_o;
  wire [3:0] n19071_o;
  wire n19072_o;
  wire n19074_o;
  wire [3:0] n19076_o;
  wire n19077_o;
  wire n19078_o;
  wire [3:0] n19079_o;
  wire n19080_o;
  wire n19081_o;
  wire [3:0] n19082_o;
  wire n19083_o;
  wire n19084_o;
  wire [3:0] n19085_o;
  wire n19086_o;
  wire n19087_o;
  wire [3:0] n19088_o;
  wire n19089_o;
  wire n19090_o;
  wire [3:0] n19091_o;
  wire n19092_o;
  wire n19093_o;
  wire [3:0] n19094_o;
  wire n19095_o;
  wire n19096_o;
  wire [7:0] n19098_o;
  wire n19099_o;
  wire n19101_o;
  wire [7:0] n19103_o;
  wire n19104_o;
  wire n19105_o;
  wire [7:0] n19106_o;
  wire n19107_o;
  wire n19108_o;
  wire [7:0] n19109_o;
  wire n19110_o;
  wire n19111_o;
  wire [15:0] n19113_o;
  wire n19114_o;
  wire n19116_o;
  wire [15:0] n19118_o;
  wire n19119_o;
  wire n19120_o;
  wire [31:0] n19122_o;
  wire n19123_o;
  wire n19125_o;
  wire [5:0] n19127_o;
  wire [3:0] n19129_o;
  wire [1:0] n19130_o;
  wire [5:0] n19131_o;
  wire n19134_o;
  wire n19135_o;
  wire [4:0] n19136_o;
  wire [5:0] n19137_o;
  wire [6:0] n19139_o;
  wire [6:0] n19141_o;
  wire [12:0] n19142_o;
  wire [12:0] n19143_o;
  wire n19146_o;
  wire [63:0] n19147_o;
  wire n19149_o;
  wire [1:0] n19150_o;
  wire [12:0] n19151_o;
  wire [63:0] n19152_o;
  wire n19153_o;
  wire n19154_o;
  localparam [63:0] n19160_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire n19163_o;
  wire n19164_o;
  wire [10:0] n19165_o;
  wire [10:0] n19167_o;
  wire [10:0] n19168_o;
  wire [10:0] n19169_o;
  wire [22:0] n19170_o;
  wire n19171_o;
  wire [28:0] n19172_o;
  wire [28:0] n19173_o;
  wire [28:0] n19174_o;
  wire n19176_o;
  wire n19179_o;
  wire n19181_o;
  wire n19182_o;
  wire [21:0] n19183_o;
  wire n19184_o;
  wire [28:0] n19185_o;
  wire [28:0] n19186_o;
  wire [28:0] n19187_o;
  wire n19189_o;
  wire [3:0] n19190_o;
  wire [28:0] n19191_o;
  reg [28:0] n19193_o;
  wire [21:0] n19194_o;
  wire [21:0] n19195_o;
  reg [21:0] n19197_o;
  wire n19198_o;
  wire n19199_o;
  reg n19201_o;
  wire [10:0] n19202_o;
  reg [10:0] n19204_o;
  wire [63:0] n19208_o;
  wire [63:0] n19209_o;
  wire n19210_o;
  wire n19212_o;
  wire [1:0] n19213_o;
  wire n19214_o;
  wire n19215_o;
  wire n19216_o;
  wire n19217_o;
  wire [4:0] n19223_o;
  wire n19225_o;
  wire n19226_o;
  wire [1:0] n19227_o;
  wire n19228_o;
  wire [2:0] n19229_o;
  wire [4:0] n19231_o;
  wire n19233_o;
  wire [1:0] n19235_o;
  wire n19236_o;
  wire [2:0] n19237_o;
  wire [4:0] n19239_o;
  wire n19241_o;
  wire n19244_o;
  wire [3:0] n19245_o;
  reg [4:0] n19247_o;
  wire [4:0] n19248_o;
  wire [4:0] n19249_o;
  wire [721:0] n19250_o;
  wire [5:0] n19251_o;
  wire n19252_o;
  wire [721:0] n19253_o;
  wire [2:0] n19254_o;
  wire n19255_o;
  wire n19256_o;
  wire [721:0] n19257_o;
  wire [4:0] n19258_o;
  wire [721:0] n19259_o;
  wire [4:0] n19260_o;
  wire [4:0] n19261_o;
  wire n19262_o;
  wire [721:0] n19263_o;
  wire [4:0] n19264_o;
  wire [4:0] n19265_o;
  wire [4:0] n19266_o;
  wire [4:0] n19267_o;
  wire n19269_o;
  wire n19270_o;
  wire n19272_o;
  wire n19273_o;
  wire [721:0] n19274_o;
  wire [3:0] n19275_o;
  wire [3:0] n19276_o;
  wire [3:0] n19277_o;
  wire n19278_o;
  wire [721:0] n19284_o;
  wire n19285_o;
  wire [721:0] n19286_o;
  wire n19287_o;
  wire n19288_o;
  wire n19289_o;
  wire n19290_o;
  wire [721:0] n19291_o;
  wire [6:0] n19292_o;
  wire n19294_o;
  wire [721:0] n19295_o;
  wire n19296_o;
  wire n19297_o;
  wire n19299_o;
  wire [9:0] n19300_o;
  wire [6:0] n19301_o;
  wire [6:0] n19302_o;
  wire n19303_o;
  wire n19304_o;
  wire n19305_o;
  wire n19306_o;
  wire n19307_o;
  wire n19308_o;
  wire n19309_o;
  wire [721:0] n19310_o;
  reg [721:0] n19318_q;
  wire [258:0] n19320_o;
  reg [18:0] n19321_q;
  wire [1:0] n19322_o;
  wire [209:0] n19323_o;
  wire [17:0] n19325_data; // mem_rd
  assign e_out_busy = n12970_o;
  assign e_out_exception = n12971_o;
  assign w_out_valid = n12973_o;
  assign w_out_interrupt = n12974_o;
  assign w_out_instr_tag = n12975_o;
  assign w_out_write_enable = n12976_o;
  assign w_out_write_reg = n12977_o;
  assign w_out_write_data = n12978_o;
  assign w_out_write_cr_enable = n12979_o;
  assign w_out_write_cr_mask = n12980_o;
  assign w_out_write_cr_data = n12981_o;
  assign w_out_intr_vec = n12982_o;
  assign w_out_srr0 = n12983_o;
  assign w_out_srr1 = n12984_o;
  /* ppc_fx_insns.vhdl:827:46  */
  assign n12968_o = {e_in_out_cr, e_in_rc, e_in_frt, e_in_frc, e_in_frb, e_in_fra, e_in_fe_mode, e_in_single, e_in_insn, e_in_itag, e_in_nia, e_in_op, e_in_valid};
  assign n12970_o = n19322_o[0];
  /* ppc_fx_insns.vhdl:766:22  */
  assign n12971_o = n19322_o[1];
  /* ppc_fx_insns.vhdl:91:18  */
  assign n12973_o = n19323_o[0];
  /* ppc_fx_insns.vhdl:91:18  */
  assign n12974_o = n19323_o[1];
  assign n12975_o = n19323_o[4:2];
  /* ppc_fx_insns.vhdl:91:18  */
  assign n12976_o = n19323_o[5];
  /* insn_helpers.vhdl:12:14  */
  assign n12977_o = n19323_o[12:6];
  /* insn_helpers.vhdl:12:14  */
  assign n12978_o = n19323_o[76:13];
  assign n12979_o = n19323_o[77];
  /* insn_helpers.vhdl:12:14  */
  assign n12980_o = n19323_o[85:78];
  /* execute1.vhdl:681:18  */
  assign n12981_o = n19323_o[117:86];
  /* insn_helpers.vhdl:22:14  */
  assign n12982_o = n19323_o[129:118];
  /* insn_helpers.vhdl:22:14  */
  assign n12983_o = n19323_o[193:130];
  assign n12984_o = n19323_o[209:194];
  /* fpu.vhdl:129:12  */
  assign r = n19318_q; // (signal)
  /* fpu.vhdl:129:15  */
  assign rin = n19310_o; // (signal)
  /* fpu.vhdl:131:12  */
  assign fp_result = n19209_o; // (signal)
  /* fpu.vhdl:132:12  */
  assign opsel_b = n16814_o; // (signal)
  /* fpu.vhdl:133:12  */
  assign opsel_r = n17513_o; // (signal)
  /* fpu.vhdl:134:12  */
  assign opsel_s = n16843_o; // (signal)
  /* fpu.vhdl:135:12  */
  assign opsel_ainv = n16847_o; // (signal)
  /* fpu.vhdl:136:12  */
  assign opsel_mask = n16852_o; // (signal)
  /* fpu.vhdl:137:12  */
  assign opsel_binv = n16857_o; // (signal)
  /* fpu.vhdl:138:12  */
  assign in_a = n18079_o; // (signal)
  /* fpu.vhdl:139:12  */
  assign in_b = n18180_o; // (signal)
  /* fpu.vhdl:140:12  */
  assign result = n18345_o; // (signal)
  /* fpu.vhdl:141:12  */
  assign carry_in = n16862_o; // (signal)
  /* fpu.vhdl:143:12  */
  assign r_hi_nz = n13500_o; // (signal)
  /* fpu.vhdl:144:12  */
  assign r_lo_nz = n13502_o; // (signal)
  /* fpu.vhdl:145:12  */
  assign s_nz = n13504_o; // (signal)
  /* fpu.vhdl:146:12  */
  assign misc_sel = n17516_o; // (signal)
  /* fpu.vhdl:147:12  */
  assign f_to_multiply = n19320_o; // (signal)
  /* fpu.vhdl:148:12  */
  assign multiply_to_f = n12991_o; // (signal)
  /* fpu.vhdl:149:12  */
  assign msel_1 = n16899_o; // (signal)
  /* fpu.vhdl:150:12  */
  assign msel_2 = n16915_o; // (signal)
  /* fpu.vhdl:151:12  */
  assign msel_add = n16925_o; // (signal)
  /* fpu.vhdl:152:12  */
  assign msel_inv = n16934_o; // (signal)
  /* fpu.vhdl:153:12  */
  assign inverse_est = n19321_q; // (signal)
  /* fpu.vhdl:535:5  */
  multiply_2 fpu_multiply_0 (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(clk),
    .m_in_valid(n12985_o),
    .m_in_data1(n12986_o),
    .m_in_data2(n12987_o),
    .m_in_addend(n12988_o),
    .m_in_is_32bit(n12989_o),
    .m_in_not_result(n12990_o),
    .m_out_valid(fpu_multiply_0_m_out_valid),
    .m_out_result(fpu_multiply_0_m_out_result),
    .m_out_overflow(fpu_multiply_0_m_out_overflow));
  /* execute1.vhdl:561:9  */
  assign n12985_o = f_to_multiply[0];
  assign n12986_o = f_to_multiply[64:1];
  /* execute1.vhdl:561:9  */
  assign n12987_o = f_to_multiply[128:65];
  assign n12988_o = f_to_multiply[256:129];
  /* execute1.vhdl:561:9  */
  assign n12989_o = f_to_multiply[257];
  assign n12990_o = f_to_multiply[258];
  /* execute1.vhdl:561:9  */
  assign n12991_o = {fpu_multiply_0_m_out_overflow, fpu_multiply_0_m_out_result, fpu_multiply_0_m_out_valid};
  /* execute1.vhdl:561:9  */
  assign n13001_o = {1'b0, 1'b0, 1'b0, 7'b0000000};
  assign n13002_o = rin[9:0];
  /* fpu.vhdl:545:13  */
  assign n13003_o = rst ? n13001_o : n13002_o;
  assign n13004_o = rin[126:10];
  /* execute1.vhdl:561:9  */
  assign n13005_o = r[126:10];
  /* fpu.vhdl:545:13  */
  assign n13006_o = rst ? n13005_o : n13004_o;
  /* execute1.vhdl:561:9  */
  assign n13007_o = rin[158:127];
  /* fpu.vhdl:545:13  */
  assign n13008_o = rst ? 32'b00000000000000000000000000000000 : n13007_o;
  /* execute1.vhdl:561:9  */
  assign n13009_o = rin[676:159];
  assign n13010_o = r[676:159];
  /* fpu.vhdl:545:13  */
  assign n13011_o = rst ? n13010_o : n13009_o;
  assign n13012_o = rin[677];
  /* fpu.vhdl:545:13  */
  assign n13013_o = rst ? 1'b0 : n13012_o;
  assign n13014_o = rin[721:678];
  /* execute1.vhdl:561:9  */
  assign n13015_o = r[721:678];
  /* fpu.vhdl:545:13  */
  assign n13016_o = rst ? n13015_o : n13014_o;
  assign n13017_o = {n13016_o, n13013_o, n13011_o, n13008_o, n13006_o, n13003_o};
  /* fpu.vhdl:565:18  */
  assign n13024_o = r[708];
  /* fpu.vhdl:566:39  */
  assign n13025_o = r[310:309];
  /* fpu.vhdl:565:13  */
  assign n13027_o = n13024_o ? n13025_o : 2'b00;
  /* fpu.vhdl:570:42  */
  assign n13028_o = r[308:301];
  /* fpu.vhdl:570:28  */
  assign n13029_o = {n13027_o, n13028_o};
  /* fpu.vhdl:571:48  */
  assign n13032_o = 10'b1111111111 - n13029_o;
  /* fpu.vhdl:571:32  */
  assign n13037_o = {1'b1, n19325_data};
  /* fpu.vhdl:575:21  */
  assign n13042_o = r[7];
  /* fpu.vhdl:576:31  */
  assign n13043_o = r[157];
  /* fpu.vhdl:578:22  */
  assign n13044_o = r[8];
  /* fpu.vhdl:578:43  */
  assign n13045_o = r[9];
  /* fpu.vhdl:578:37  */
  assign n13046_o = ~n13045_o;
  /* fpu.vhdl:578:33  */
  assign n13047_o = n13044_o & n13046_o;
  /* fpu.vhdl:579:26  */
  assign n13048_o = r[115:113];
  /* fpu.vhdl:580:29  */
  assign n13049_o = r[677];
  /* fpu.vhdl:581:26  */
  assign n13050_o = r[122:116];
  /* fpu.vhdl:583:32  */
  assign n13051_o = r[8];
  /* fpu.vhdl:583:50  */
  assign n13052_o = r[124];
  /* fpu.vhdl:583:58  */
  assign n13053_o = r[125];
  /* fpu.vhdl:583:53  */
  assign n13054_o = n13052_o | n13053_o;
  /* fpu.vhdl:583:43  */
  assign n13055_o = n13051_o & n13054_o;
  /* fpu.vhdl:584:30  */
  assign n13056_o = r[690:683];
  /* fpu.vhdl:585:30  */
  assign n13057_o = r[682:679];
  /* fpu.vhdl:585:44  */
  assign n13058_o = r[682:679];
  /* fpu.vhdl:585:40  */
  assign n13059_o = {n13057_o, n13058_o};
  /* fpu.vhdl:585:58  */
  assign n13060_o = r[682:679];
  /* fpu.vhdl:585:54  */
  assign n13061_o = {n13059_o, n13060_o};
  /* fpu.vhdl:585:72  */
  assign n13062_o = r[682:679];
  /* fpu.vhdl:585:68  */
  assign n13063_o = {n13061_o, n13062_o};
  /* fpu.vhdl:586:30  */
  assign n13064_o = r[682:679];
  /* fpu.vhdl:585:82  */
  assign n13065_o = {n13063_o, n13064_o};
  /* fpu.vhdl:586:44  */
  assign n13066_o = r[682:679];
  /* fpu.vhdl:586:40  */
  assign n13067_o = {n13065_o, n13066_o};
  /* fpu.vhdl:586:58  */
  assign n13068_o = r[682:679];
  /* fpu.vhdl:586:54  */
  assign n13069_o = {n13067_o, n13068_o};
  /* fpu.vhdl:586:72  */
  assign n13070_o = r[682:679];
  /* fpu.vhdl:586:68  */
  assign n13071_o = {n13069_o, n13070_o};
  /* fpu.vhdl:587:26  */
  assign n13072_o = r[9];
  /* fpu.vhdl:589:21  */
  assign n13074_o = r[112:49];
  /* fpu.vhdl:590:31  */
  assign n13075_o = r[10];
  /* fpu.vhdl:590:55  */
  assign n13076_o = r[10];
  /* fpu.vhdl:590:49  */
  assign n13077_o = ~n13076_o;
  assign n13092_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* execute1.vhdl:451:18  */
  assign n13093_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n13094_o = {1'b0, 1'b0, 1'b0, n13077_o};
  /* execute1.vhdl:450:18  */
  assign n13095_o = {n13075_o, 1'b0, 1'b0, 1'b0};
  assign n13096_o = {n13092_o, n13093_o, n13094_o, n13095_o};
  assign n13151_o = r[6:0];
  /* fpu.vhdl:650:17  */
  assign n13152_o = n12968_o[0];
  /* fpu.vhdl:651:28  */
  assign n13153_o = n12968_o[105:74];
  /* fpu.vhdl:652:27  */
  assign n13154_o = n12968_o[70:7];
  /* fpu.vhdl:653:26  */
  assign n13155_o = n12968_o[6:1];
  /* fpu.vhdl:654:33  */
  assign n13156_o = n12968_o[73:71];
  /* fpu.vhdl:655:35  */
  assign n13157_o = n12968_o[108:107];
  /* fpu.vhdl:655:26  */
  assign n13158_o = |(n13157_o);
  /* fpu.vhdl:656:32  */
  assign n13159_o = n12968_o[307:301];
  /* fpu.vhdl:657:35  */
  assign n13160_o = n12968_o[106];
  /* fpu.vhdl:658:32  */
  assign n13161_o = n12968_o[106];
  /* fpu.vhdl:660:26  */
  assign n13163_o = n12968_o[308];
  /* fpu.vhdl:661:30  */
  assign n13164_o = n12968_o[309];
  /* fpu.vhdl:662:21  */
  assign n13165_o = n12968_o[309];
  /* fpu.vhdl:662:28  */
  assign n13166_o = ~n13165_o;
  /* fpu.vhdl:665:74  */
  assign n13171_o = n12968_o[105:74];
  /* insn_helpers.vhdl:136:23  */
  assign n13176_o = n13171_o[25:23];
  /* crhelpers.vhdl:36:13  */
  assign n13184_o = n13176_o == 3'b000;
  /* crhelpers.vhdl:38:13  */
  assign n13187_o = n13176_o == 3'b001;
  /* crhelpers.vhdl:40:13  */
  assign n13190_o = n13176_o == 3'b010;
  /* crhelpers.vhdl:42:13  */
  assign n13193_o = n13176_o == 3'b011;
  /* crhelpers.vhdl:44:13  */
  assign n13196_o = n13176_o == 3'b100;
  /* crhelpers.vhdl:46:13  */
  assign n13199_o = n13176_o == 3'b101;
  /* crhelpers.vhdl:48:13  */
  assign n13202_o = n13176_o == 3'b110;
  /* crhelpers.vhdl:50:13  */
  assign n13205_o = n13176_o == 3'b111;
  assign n13207_o = {n13205_o, n13202_o, n13199_o, n13196_o, n13193_o, n13190_o, n13187_o, n13184_o};
  /* crhelpers.vhdl:35:9  */
  always @*
    case (n13207_o)
      8'b10000000: n13208_o = 8'b00000001;
      8'b01000000: n13208_o = 8'b00000010;
      8'b00100000: n13208_o = 8'b00000100;
      8'b00010000: n13208_o = 8'b00001000;
      8'b00001000: n13208_o = 8'b00010000;
      8'b00000100: n13208_o = 8'b00100000;
      8'b00000010: n13208_o = 8'b01000000;
      8'b00000001: n13208_o = 8'b10000000;
      default: n13208_o = 8'b00000000;
    endcase
  /* fpu.vhdl:662:13  */
  assign n13209_o = n13166_o ? 8'b01000000 : n13208_o;
  /* fpu.vhdl:668:21  */
  assign n13210_o = n12968_o[6:1];
  /* fpu.vhdl:668:24  */
  assign n13212_o = n13210_o == 6'b011010;
  /* fpu.vhdl:668:13  */
  assign n13215_o = n13212_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:674:42  */
  assign n13220_o = r[128:127];
  /* fpu.vhdl:674:33  */
  assign n13222_o = {1'b0, n13220_o};
  /* fpu.vhdl:681:36  */
  assign n13229_o = n12968_o[172:109];
  /* fpu.vhdl:417:26  */
  assign n13239_o = n13229_o[63];
  /* fpu.vhdl:418:26  */
  assign n13243_o = n13229_o[62:52];
  /* fpu.vhdl:418:19  */
  assign n13244_o = |(n13243_o);
  /* fpu.vhdl:419:27  */
  assign n13246_o = n13229_o[62:52];
  /* fpu.vhdl:419:19  */
  assign n13247_o = &(n13246_o);
  /* fpu.vhdl:420:27  */
  assign n13249_o = n13229_o[51:0];
  /* fpu.vhdl:420:20  */
  assign n13250_o = |(n13249_o);
  /* fpu.vhdl:421:19  */
  assign n13252_o = ~n13215_o;
  /* fpu.vhdl:422:53  */
  assign n13253_o = n13229_o[62:52];
  /* fpu.vhdl:422:34  */
  assign n13254_o = {2'b0, n13253_o};  //  uext
  /* fpu.vhdl:422:81  */
  assign n13256_o = n13254_o - 13'b0001111111111;
  /* fpu.vhdl:423:23  */
  assign n13257_o = ~n13244_o;
  /* fpu.vhdl:423:13  */
  assign n13259_o = n13257_o ? 13'b1110000000010 : n13256_o;
  /* fpu.vhdl:426:39  */
  assign n13261_o = {9'b000000000, n13244_o};
  /* fpu.vhdl:426:53  */
  assign n13262_o = n13229_o[51:0];
  /* fpu.vhdl:426:48  */
  assign n13263_o = {n13261_o, n13262_o};
  /* fpu.vhdl:426:67  */
  assign n13265_o = {n13263_o, 2'b00};
  /* fpu.vhdl:427:27  */
  assign n13266_o = {n13247_o, n13244_o};
  /* fpu.vhdl:427:36  */
  assign n13267_o = {n13266_o, n13250_o};
  /* fpu.vhdl:429:17  */
  assign n13270_o = n13267_o == 3'b000;
  /* fpu.vhdl:430:17  */
  assign n13273_o = n13267_o == 3'b001;
  /* fpu.vhdl:431:17  */
  assign n13276_o = n13267_o == 3'b010;
  /* fpu.vhdl:432:17  */
  assign n13279_o = n13267_o == 3'b011;
  /* fpu.vhdl:433:17  */
  assign n13282_o = n13267_o == 3'b110;
  assign n13284_o = {n13282_o, n13279_o, n13276_o, n13273_o, n13270_o};
  /* fpu.vhdl:428:13  */
  always @*
    case (n13284_o)
      5'b10000: n13285_o = 2'b10;
      5'b01000: n13285_o = 2'b01;
      5'b00100: n13285_o = 2'b01;
      5'b00010: n13285_o = 2'b01;
      5'b00001: n13285_o = 2'b00;
      default: n13285_o = 2'b11;
    endcase
  /* fpu.vhdl:439:20  */
  assign n13287_o = n13229_o[63];
  /* fpu.vhdl:439:25  */
  assign n13288_o = n13287_o | n13244_o;
  /* fpu.vhdl:439:35  */
  assign n13289_o = n13288_o | n13250_o;
  /* fpu.vhdl:439:13  */
  assign n13292_o = n13289_o ? 2'b01 : 2'b00;
  assign n13293_o = {n13229_o, 13'b0000000000000};
  assign n13294_o = {n13265_o, n13259_o};
  /* fpu.vhdl:421:9  */
  assign n13295_o = n13252_o ? n13285_o : n13292_o;
  /* fpu.vhdl:421:9  */
  assign n13296_o = n13252_o ? n13294_o : n13293_o;
  assign n13300_o = {n13296_o, n13239_o, n13295_o};
  /* fpu.vhdl:682:36  */
  assign n13302_o = n12968_o[236:173];
  /* fpu.vhdl:417:26  */
  assign n13312_o = n13302_o[63];
  /* fpu.vhdl:418:26  */
  assign n13316_o = n13302_o[62:52];
  /* fpu.vhdl:418:19  */
  assign n13317_o = |(n13316_o);
  /* fpu.vhdl:419:27  */
  assign n13319_o = n13302_o[62:52];
  /* fpu.vhdl:419:19  */
  assign n13320_o = &(n13319_o);
  /* fpu.vhdl:420:27  */
  assign n13322_o = n13302_o[51:0];
  /* fpu.vhdl:420:20  */
  assign n13323_o = |(n13322_o);
  /* fpu.vhdl:421:19  */
  assign n13325_o = ~n13215_o;
  /* fpu.vhdl:422:53  */
  assign n13326_o = n13302_o[62:52];
  /* fpu.vhdl:422:34  */
  assign n13327_o = {2'b0, n13326_o};  //  uext
  /* fpu.vhdl:422:81  */
  assign n13329_o = n13327_o - 13'b0001111111111;
  /* fpu.vhdl:423:23  */
  assign n13330_o = ~n13317_o;
  /* fpu.vhdl:423:13  */
  assign n13332_o = n13330_o ? 13'b1110000000010 : n13329_o;
  /* fpu.vhdl:426:39  */
  assign n13334_o = {9'b000000000, n13317_o};
  /* fpu.vhdl:426:53  */
  assign n13335_o = n13302_o[51:0];
  /* fpu.vhdl:426:48  */
  assign n13336_o = {n13334_o, n13335_o};
  /* fpu.vhdl:426:67  */
  assign n13338_o = {n13336_o, 2'b00};
  /* fpu.vhdl:427:27  */
  assign n13339_o = {n13320_o, n13317_o};
  /* fpu.vhdl:427:36  */
  assign n13340_o = {n13339_o, n13323_o};
  /* fpu.vhdl:429:17  */
  assign n13343_o = n13340_o == 3'b000;
  /* fpu.vhdl:430:17  */
  assign n13346_o = n13340_o == 3'b001;
  /* fpu.vhdl:431:17  */
  assign n13349_o = n13340_o == 3'b010;
  /* fpu.vhdl:432:17  */
  assign n13352_o = n13340_o == 3'b011;
  /* fpu.vhdl:433:17  */
  assign n13355_o = n13340_o == 3'b110;
  assign n13357_o = {n13355_o, n13352_o, n13349_o, n13346_o, n13343_o};
  /* fpu.vhdl:428:13  */
  always @*
    case (n13357_o)
      5'b10000: n13358_o = 2'b10;
      5'b01000: n13358_o = 2'b01;
      5'b00100: n13358_o = 2'b01;
      5'b00010: n13358_o = 2'b01;
      5'b00001: n13358_o = 2'b00;
      default: n13358_o = 2'b11;
    endcase
  /* fpu.vhdl:439:20  */
  assign n13360_o = n13302_o[63];
  /* fpu.vhdl:439:25  */
  assign n13361_o = n13360_o | n13317_o;
  /* fpu.vhdl:439:35  */
  assign n13362_o = n13361_o | n13323_o;
  /* fpu.vhdl:439:13  */
  assign n13365_o = n13362_o ? 2'b01 : 2'b00;
  assign n13366_o = {n13302_o, 13'b0000000000000};
  assign n13367_o = {n13338_o, n13332_o};
  /* fpu.vhdl:421:9  */
  assign n13368_o = n13325_o ? n13358_o : n13365_o;
  /* fpu.vhdl:421:9  */
  assign n13369_o = n13325_o ? n13367_o : n13366_o;
  assign n13373_o = {n13369_o, n13312_o, n13368_o};
  /* fpu.vhdl:683:36  */
  assign n13375_o = n12968_o[300:237];
  /* fpu.vhdl:417:26  */
  assign n13385_o = n13375_o[63];
  /* fpu.vhdl:418:26  */
  assign n13389_o = n13375_o[62:52];
  /* fpu.vhdl:418:19  */
  assign n13390_o = |(n13389_o);
  /* fpu.vhdl:419:27  */
  assign n13392_o = n13375_o[62:52];
  /* fpu.vhdl:419:19  */
  assign n13393_o = &(n13392_o);
  /* fpu.vhdl:420:27  */
  assign n13395_o = n13375_o[51:0];
  /* fpu.vhdl:420:20  */
  assign n13396_o = |(n13395_o);
  /* fpu.vhdl:421:19  */
  assign n13398_o = ~n13215_o;
  /* fpu.vhdl:422:53  */
  assign n13399_o = n13375_o[62:52];
  /* fpu.vhdl:422:34  */
  assign n13400_o = {2'b0, n13399_o};  //  uext
  /* fpu.vhdl:422:81  */
  assign n13402_o = n13400_o - 13'b0001111111111;
  /* fpu.vhdl:423:23  */
  assign n13403_o = ~n13390_o;
  /* fpu.vhdl:423:13  */
  assign n13405_o = n13403_o ? 13'b1110000000010 : n13402_o;
  /* fpu.vhdl:426:39  */
  assign n13407_o = {9'b000000000, n13390_o};
  /* fpu.vhdl:426:53  */
  assign n13408_o = n13375_o[51:0];
  /* fpu.vhdl:426:48  */
  assign n13409_o = {n13407_o, n13408_o};
  /* fpu.vhdl:426:67  */
  assign n13411_o = {n13409_o, 2'b00};
  /* fpu.vhdl:427:27  */
  assign n13412_o = {n13393_o, n13390_o};
  /* fpu.vhdl:427:36  */
  assign n13413_o = {n13412_o, n13396_o};
  /* fpu.vhdl:429:17  */
  assign n13416_o = n13413_o == 3'b000;
  /* fpu.vhdl:430:17  */
  assign n13419_o = n13413_o == 3'b001;
  /* fpu.vhdl:431:17  */
  assign n13422_o = n13413_o == 3'b010;
  /* fpu.vhdl:432:17  */
  assign n13425_o = n13413_o == 3'b011;
  /* fpu.vhdl:433:17  */
  assign n13428_o = n13413_o == 3'b110;
  assign n13430_o = {n13428_o, n13425_o, n13422_o, n13419_o, n13416_o};
  /* fpu.vhdl:428:13  */
  always @*
    case (n13430_o)
      5'b10000: n13431_o = 2'b10;
      5'b01000: n13431_o = 2'b01;
      5'b00100: n13431_o = 2'b01;
      5'b00010: n13431_o = 2'b01;
      5'b00001: n13431_o = 2'b00;
      default: n13431_o = 2'b11;
    endcase
  /* fpu.vhdl:439:20  */
  assign n13433_o = n13375_o[63];
  /* fpu.vhdl:439:25  */
  assign n13434_o = n13433_o | n13390_o;
  /* fpu.vhdl:439:35  */
  assign n13435_o = n13434_o | n13396_o;
  /* fpu.vhdl:439:13  */
  assign n13438_o = n13435_o ? 2'b01 : 2'b00;
  assign n13439_o = {n13375_o, 13'b0000000000000};
  assign n13440_o = {n13411_o, n13405_o};
  /* fpu.vhdl:421:9  */
  assign n13441_o = n13398_o ? n13431_o : n13438_o;
  /* fpu.vhdl:421:9  */
  assign n13442_o = n13398_o ? n13440_o : n13439_o;
  assign n13446_o = {n13442_o, n13385_o, n13441_o};
  /* fpu.vhdl:689:21  */
  assign n13448_o = n13300_o[15:3];
  /* fpu.vhdl:689:37  */
  assign n13449_o = n13373_o[15:3];
  /* fpu.vhdl:689:30  */
  assign n13450_o = $signed(n13448_o) > $signed(n13449_o);
  /* fpu.vhdl:689:13  */
  assign n13452_o = n13450_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:693:22  */
  assign n13454_o = n13300_o[15:3];
  /* fpu.vhdl:693:38  */
  assign n13455_o = n13446_o[15:3];
  /* fpu.vhdl:693:31  */
  assign n13456_o = n13454_o + n13455_o;
  /* fpu.vhdl:693:47  */
  assign n13458_o = n13456_o + 13'b0000000000001;
  /* fpu.vhdl:693:60  */
  assign n13459_o = n13373_o[15:3];
  /* fpu.vhdl:693:52  */
  assign n13460_o = $signed(n13458_o) >= $signed(n13459_o);
  /* fpu.vhdl:693:13  */
  assign n13462_o = n13460_o ? 1'b1 : 1'b0;
  assign n13463_o = {n13160_o, n13164_o, n13163_o, n13158_o, n13159_o, n13156_o, n13154_o, n13153_o, n13155_o};
  assign n13464_o = {n13446_o, n13373_o, n13300_o};
  assign n13465_o = {1'b0, 1'b0, 1'b0, n13462_o, n13452_o, 1'b0, n13222_o, 1'b0, 1'b0, 1'b1};
  assign n13466_o = r[126:11];
  /* fpu.vhdl:650:9  */
  assign n13467_o = n13152_o ? n13463_o : n13466_o;
  assign n13468_o = r[398:159];
  /* fpu.vhdl:650:9  */
  assign n13469_o = n13152_o ? n13464_o : n13468_o;
  assign n13470_o = r[678];
  /* fpu.vhdl:650:9  */
  assign n13471_o = n13152_o ? 1'b0 : n13470_o;
  assign n13472_o = r[690:683];
  /* fpu.vhdl:650:9  */
  assign n13473_o = n13152_o ? n13209_o : n13472_o;
  assign n13474_o = r[708:697];
  /* fpu.vhdl:650:9  */
  assign n13475_o = n13152_o ? n13465_o : n13474_o;
  assign n13476_o = r[713:712];
  /* fpu.vhdl:650:9  */
  assign n13477_o = n13152_o ? 2'b00 : n13476_o;
  assign n13478_o = r[721];
  /* fpu.vhdl:650:9  */
  assign n13479_o = n13152_o ? n13161_o : n13478_o;
  assign n13483_o = r[158:127];
  assign n13487_o = r[682:679];
  /* fpu.vhdl:650:9  */
  assign n13497_o = n13152_o ? n13215_o : 1'b0;
  /* fpu.vhdl:698:27  */
  assign n13499_o = r[454:430];
  /* fpu.vhdl:698:20  */
  assign n13500_o = |(n13499_o);
  /* fpu.vhdl:699:27  */
  assign n13501_o = r[429:401];
  /* fpu.vhdl:699:20  */
  assign n13502_o = |(n13501_o);
  /* fpu.vhdl:700:23  */
  assign n13503_o = r[518:463];
  /* fpu.vhdl:700:17  */
  assign n13504_o = |(n13503_o);
  /* fpu.vhdl:702:14  */
  assign n13505_o = r[126];
  /* fpu.vhdl:702:26  */
  assign n13506_o = ~n13505_o;
  /* fpu.vhdl:703:29  */
  assign n13507_o = r[713];
  /* fpu.vhdl:703:33  */
  assign n13508_o = ~n13507_o;
  /* fpu.vhdl:703:13  */
  assign n13511_o = n13508_o ? 13'b0001111111111 : 13'b0001111111100;
  /* fpu.vhdl:708:29  */
  assign n13512_o = r[712];
  /* fpu.vhdl:708:33  */
  assign n13513_o = ~n13512_o;
  /* fpu.vhdl:708:13  */
  assign n13516_o = n13513_o ? 13'b1110000000010 : 13'b1110000000011;
  /* fpu.vhdl:702:9  */
  assign n13518_o = n13506_o ? n13516_o : 13'b1111110000010;
  /* fpu.vhdl:702:9  */
  assign n13520_o = n13506_o ? n13511_o : 13'b0000001111111;
  /* fpu.vhdl:702:9  */
  assign n13523_o = n13506_o ? 13'b0011000000000 : 13'b0000011000000;
  /* fpu.vhdl:719:22  */
  assign n13524_o = r[663:651];
  /* fpu.vhdl:719:37  */
  assign n13525_o = r[676:664];
  /* fpu.vhdl:719:33  */
  assign n13526_o = n13524_o - n13525_o;
  /* fpu.vhdl:722:20  */
  assign n13527_o = $signed(n13526_o) < $signed(n13518_o);
  /* fpu.vhdl:722:9  */
  assign n13530_o = n13527_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:725:20  */
  assign n13532_o = $signed(n13526_o) > $signed(n13520_o);
  /* fpu.vhdl:725:9  */
  assign n13535_o = n13532_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:730:25  */
  assign n13537_o = r[577:524];
  /* fpu.vhdl:730:18  */
  assign n13538_o = |(n13537_o);
  /* fpu.vhdl:732:15  */
  assign n13539_o = r[579:524];
  /* fpu.vhdl:732:43  */
  assign n13540_o = r[310:255];
  /* fpu.vhdl:732:29  */
  assign n13541_o = n13539_o == n13540_o;
  /* fpu.vhdl:732:9  */
  assign n13544_o = n13541_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:736:24  */
  assign n13546_o = r[579:524];
  /* fpu.vhdl:736:62  */
  assign n13547_o = r[310:255];
  /* fpu.vhdl:736:39  */
  assign n13548_o = $unsigned(n13546_o) < $unsigned(n13547_o);
  /* fpu.vhdl:736:9  */
  assign n13551_o = n13548_o ? 1'b1 : 1'b0;
  assign n13556_o = r[10:9];
  assign n13558_o = r[695:691];
  assign n13560_o = r[663:399];
  assign n13562_o = r[711:710];
  assign n13564_o = r[720:716];
  /* fpu.vhdl:776:16  */
  assign n13567_o = r[6:0];
  /* fpu.vhdl:783:25  */
  assign n13573_o = n12968_o[0];
  /* fpu.vhdl:784:35  */
  assign n13574_o = n12968_o[79:75];
  /* fpu.vhdl:786:41  */
  assign n13575_o = n12968_o[82];
  /* fpu.vhdl:787:45  */
  assign n13576_o = n12968_o[80];
  /* fpu.vhdl:787:49  */
  assign n13577_o = ~n13576_o;
  /* fpu.vhdl:787:33  */
  assign n13580_o = n13577_o ? 7'b0001001 : 7'b0001010;
  /* fpu.vhdl:792:44  */
  assign n13581_o = n12968_o[81];
  /* fpu.vhdl:792:29  */
  assign n13585_o = n13581_o ? 7'b0000001 : 7'b0001000;
  /* fpu.vhdl:792:29  */
  assign n13586_o = n13581_o ? 2'b00 : 2'b10;
  /* fpu.vhdl:786:29  */
  assign n13587_o = n13575_o ? n13580_o : n13585_o;
  /* fpu.vhdl:786:29  */
  assign n13588_o = n13575_o ? 2'b00 : n13586_o;
  /* fpu.vhdl:785:25  */
  assign n13590_o = n13574_o == 5'b00000;
  /* fpu.vhdl:799:41  */
  assign n13591_o = n12968_o[84];
  /* fpu.vhdl:799:46  */
  assign n13592_o = ~n13591_o;
  /* fpu.vhdl:800:45  */
  assign n13593_o = n12968_o[82];
  /* fpu.vhdl:800:49  */
  assign n13594_o = ~n13593_o;
  /* fpu.vhdl:800:33  */
  assign n13597_o = n13594_o ? 7'b0000010 : 7'b0000011;
  /* fpu.vhdl:799:29  */
  assign n13599_o = n13592_o ? n13597_o : 7'b0000111;
  /* fpu.vhdl:798:25  */
  assign n13601_o = n13574_o == 5'b00110;
  /* fpu.vhdl:809:41  */
  assign n13602_o = n12968_o[82];
  /* fpu.vhdl:809:45  */
  assign n13603_o = ~n13602_o;
  /* fpu.vhdl:809:29  */
  assign n13606_o = n13603_o ? 7'b0000100 : 7'b0000101;
  /* fpu.vhdl:808:25  */
  assign n13608_o = n13574_o == 5'b00111;
  /* fpu.vhdl:816:41  */
  assign n13610_o = n12968_o[83:82];
  /* fpu.vhdl:816:54  */
  assign n13612_o = n13610_o != 2'b11;
  /* fpu.vhdl:816:29  */
  assign n13615_o = n13612_o ? 7'b0000110 : 7'b0001110;
  /* fpu.vhdl:814:25  */
  assign n13617_o = n13574_o == 5'b01000;
  /* fpu.vhdl:821:25  */
  assign n13621_o = n13574_o == 5'b01100;
  /* fpu.vhdl:826:29  */
  assign n13625_o = n13497_o ? 7'b0001011 : 7'b0001100;
  /* fpu.vhdl:824:25  */
  assign n13627_o = n13574_o == 5'b01110;
  /* fpu.vhdl:832:25  */
  assign n13632_o = n13574_o == 5'b01111;
  assign n13634_o = {n13479_o, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, n13477_o, n13562_o, 1'b0, n13475_o, 1'b0, n13558_o, n13473_o, n13487_o, n13471_o, 1'b0, 13'b0000000000000, n13560_o, n13469_o, n13483_o, n13467_o, n13556_o, 1'b0, 1'b0, n13151_o};
  /* fpu.vhdl:838:44  */
  assign n13635_o = n13634_o[309];
  /* fpu.vhdl:838:49  */
  assign n13636_o = ~n13635_o;
  assign n13637_o = {n13479_o, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, n13477_o, n13562_o, 1'b0, n13475_o, 1'b0, n13558_o, n13473_o, n13487_o, n13471_o, 1'b0, 13'b0000000000000, n13560_o, n13469_o, n13483_o, n13467_o, n13556_o, 1'b0, 1'b0, n13151_o};
  /* fpu.vhdl:838:71  */
  assign n13638_o = n13637_o[229];
  /* fpu.vhdl:838:55  */
  assign n13639_o = n13636_o & n13638_o;
  /* fpu.vhdl:838:29  */
  assign n13641_o = n13639_o ? 2'b10 : 2'b01;
  /* fpu.vhdl:836:25  */
  assign n13644_o = n13574_o == 5'b10010;
  /* fpu.vhdl:842:25  */
  assign n13648_o = n13574_o == 5'b10100;
  /* fpu.vhdl:842:38  */
  assign n13650_o = n13574_o == 5'b10101;
  /* fpu.vhdl:842:38  */
  assign n13651_o = n13648_o | n13650_o;
  /* fpu.vhdl:845:25  */
  assign n13656_o = n13574_o == 5'b10110;
  /* fpu.vhdl:849:25  */
  assign n13659_o = n13574_o == 5'b10111;
  /* fpu.vhdl:851:25  */
  assign n13663_o = n13574_o == 5'b11000;
  assign n13666_o = n13465_o[9:0];
  assign n13667_o = r[706:697];
  /* fpu.vhdl:650:9  */
  assign n13668_o = n13152_o ? n13666_o : n13667_o;
  assign n13669_o = n13465_o[11];
  assign n13670_o = r[708];
  /* fpu.vhdl:650:9  */
  assign n13671_o = n13152_o ? n13669_o : n13670_o;
  assign n13672_o = {n13479_o, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, n13477_o, n13562_o, 1'b0, n13671_o, 1'b1, n13668_o, 1'b0, n13558_o, n13473_o, n13487_o, n13471_o, 1'b0, 13'b0000000000000, n13560_o, n13469_o, n13483_o, n13467_o, n13556_o, 1'b0, 1'b0, n13151_o};
  /* fpu.vhdl:857:44  */
  assign n13673_o = n13672_o[389];
  /* fpu.vhdl:857:49  */
  assign n13674_o = ~n13673_o;
  assign n13675_o = n13465_o[9:0];
  assign n13676_o = r[706:697];
  /* fpu.vhdl:650:9  */
  assign n13677_o = n13152_o ? n13675_o : n13676_o;
  assign n13678_o = n13465_o[11];
  assign n13679_o = r[708];
  /* fpu.vhdl:650:9  */
  assign n13680_o = n13152_o ? n13678_o : n13679_o;
  assign n13681_o = {n13479_o, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 2'b01, n13477_o, n13562_o, 1'b0, n13680_o, 1'b1, n13677_o, 1'b0, n13558_o, n13473_o, n13487_o, n13471_o, 1'b0, 13'b0000000000000, n13560_o, n13469_o, n13483_o, n13467_o, n13556_o, 1'b0, 1'b0, n13151_o};
  /* fpu.vhdl:857:71  */
  assign n13682_o = n13681_o[229];
  /* fpu.vhdl:857:55  */
  assign n13683_o = n13674_o & n13682_o;
  /* fpu.vhdl:857:29  */
  assign n13685_o = n13683_o ? 2'b11 : 2'b01;
  /* fpu.vhdl:854:25  */
  assign n13688_o = n13574_o == 5'b11001;
  /* fpu.vhdl:861:25  */
  assign n13693_o = n13574_o == 5'b11010;
  assign n13694_o = {n13479_o, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, n13477_o, n13562_o, 1'b0, n13475_o, 1'b0, n13558_o, n13473_o, n13487_o, n13471_o, 1'b0, 13'b0000000000000, n13560_o, n13469_o, n13483_o, n13467_o, n13556_o, 1'b0, 1'b0, n13151_o};
  /* fpu.vhdl:866:44  */
  assign n13695_o = n13694_o[229];
  /* fpu.vhdl:866:49  */
  assign n13696_o = ~n13695_o;
  assign n13698_o = {n13479_o, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 2'b00, n13477_o, n13562_o, 1'b0, n13475_o, 1'b0, n13558_o, n13473_o, n13487_o, n13471_o, 1'b0, 13'b0000000000000, n13560_o, n13469_o, n13483_o, n13467_o, n13556_o, 1'b0, 1'b0, n13151_o};
  /* fpu.vhdl:868:47  */
  assign n13699_o = n13698_o[389];
  /* fpu.vhdl:868:52  */
  assign n13700_o = ~n13699_o;
  /* fpu.vhdl:868:29  */
  assign n13703_o = n13700_o ? 2'b11 : 2'b10;
  /* fpu.vhdl:866:29  */
  assign n13704_o = n13696_o ? 2'b01 : n13703_o;
  /* fpu.vhdl:865:25  */
  assign n13707_o = n13574_o == 5'b11100;
  /* fpu.vhdl:865:38  */
  assign n13709_o = n13574_o == 5'b11101;
  /* fpu.vhdl:865:38  */
  assign n13710_o = n13707_o | n13709_o;
  /* fpu.vhdl:865:48  */
  assign n13712_o = n13574_o == 5'b11110;
  /* fpu.vhdl:865:48  */
  assign n13713_o = n13710_o | n13712_o;
  /* fpu.vhdl:865:58  */
  assign n13715_o = n13574_o == 5'b11111;
  /* fpu.vhdl:865:58  */
  assign n13716_o = n13713_o | n13715_o;
  assign n13717_o = {n13716_o, n13693_o, n13688_o, n13663_o, n13659_o, n13656_o, n13651_o, n13644_o, n13632_o, n13627_o, n13621_o, n13617_o, n13608_o, n13601_o, n13590_o};
  /* fpu.vhdl:784:21  */
  always @*
    case (n13717_o)
      15'b100000000000000: n13718_o = 7'b0010011;
      15'b010000000000000: n13718_o = 7'b0010101;
      15'b001000000000000: n13718_o = 7'b0010000;
      15'b000100000000000: n13718_o = 7'b0010100;
      15'b000010000000000: n13718_o = 7'b0010110;
      15'b000001000000000: n13718_o = 7'b0010010;
      15'b000000100000000: n13718_o = 7'b0001111;
      15'b000000010000000: n13718_o = 7'b0010001;
      15'b000000001000000: n13718_o = 7'b0001100;
      15'b000000000100000: n13718_o = n13625_o;
      15'b000000000010000: n13718_o = 7'b0001101;
      15'b000000000001000: n13718_o = n13615_o;
      15'b000000000000100: n13718_o = n13606_o;
      15'b000000000000010: n13718_o = n13599_o;
      15'b000000000000001: n13718_o = n13587_o;
      default: n13718_o = n13151_o;
    endcase
  assign n13719_o = n13465_o[5:3];
  assign n13720_o = r[702:700];
  /* fpu.vhdl:650:9  */
  assign n13721_o = n13152_o ? n13719_o : n13720_o;
  /* fpu.vhdl:784:21  */
  always @*
    case (n13717_o)
      15'b100000000000000: n13722_o = n13721_o;
      15'b010000000000000: n13722_o = n13721_o;
      15'b001000000000000: n13722_o = n13721_o;
      15'b000100000000000: n13722_o = n13721_o;
      15'b000010000000000: n13722_o = n13721_o;
      15'b000001000000000: n13722_o = n13721_o;
      15'b000000100000000: n13722_o = n13721_o;
      15'b000000010000000: n13722_o = n13721_o;
      15'b000000001000000: n13722_o = 3'b001;
      15'b000000000100000: n13722_o = n13721_o;
      15'b000000000010000: n13722_o = n13721_o;
      15'b000000000001000: n13722_o = n13721_o;
      15'b000000000000100: n13722_o = n13721_o;
      15'b000000000000010: n13722_o = n13721_o;
      15'b000000000000001: n13722_o = n13721_o;
      default: n13722_o = n13721_o;
    endcase
  assign n13723_o = n13465_o[10];
  assign n13724_o = r[707];
  /* fpu.vhdl:650:9  */
  assign n13725_o = n13152_o ? n13723_o : n13724_o;
  /* fpu.vhdl:784:21  */
  always @*
    case (n13717_o)
      15'b100000000000000: n13726_o = n13725_o;
      15'b010000000000000: n13726_o = n13725_o;
      15'b001000000000000: n13726_o = 1'b1;
      15'b000100000000000: n13726_o = n13725_o;
      15'b000010000000000: n13726_o = n13725_o;
      15'b000001000000000: n13726_o = n13725_o;
      15'b000000100000000: n13726_o = n13725_o;
      15'b000000010000000: n13726_o = n13725_o;
      15'b000000001000000: n13726_o = n13725_o;
      15'b000000000100000: n13726_o = n13725_o;
      15'b000000000010000: n13726_o = n13725_o;
      15'b000000000001000: n13726_o = n13725_o;
      15'b000000000000100: n13726_o = n13725_o;
      15'b000000000000010: n13726_o = n13725_o;
      15'b000000000000001: n13726_o = n13725_o;
      default: n13726_o = n13725_o;
    endcase
  assign n13727_o = n13465_o[11];
  assign n13728_o = r[708];
  /* fpu.vhdl:650:9  */
  assign n13729_o = n13152_o ? n13727_o : n13728_o;
  /* fpu.vhdl:784:21  */
  always @*
    case (n13717_o)
      15'b100000000000000: n13730_o = n13729_o;
      15'b010000000000000: n13730_o = 1'b1;
      15'b001000000000000: n13730_o = n13729_o;
      15'b000100000000000: n13730_o = n13729_o;
      15'b000010000000000: n13730_o = n13729_o;
      15'b000001000000000: n13730_o = 1'b1;
      15'b000000100000000: n13730_o = n13729_o;
      15'b000000010000000: n13730_o = n13729_o;
      15'b000000001000000: n13730_o = n13729_o;
      15'b000000000100000: n13730_o = n13729_o;
      15'b000000000010000: n13730_o = n13729_o;
      15'b000000000001000: n13730_o = n13729_o;
      15'b000000000000100: n13730_o = n13729_o;
      15'b000000000000010: n13730_o = n13729_o;
      15'b000000000000001: n13730_o = n13729_o;
      default: n13730_o = n13729_o;
    endcase
  /* fpu.vhdl:784:21  */
  always @*
    case (n13717_o)
      15'b100000000000000: n13731_o = n13704_o;
      15'b010000000000000: n13731_o = 2'b10;
      15'b001000000000000: n13731_o = n13685_o;
      15'b000100000000000: n13731_o = 2'b10;
      15'b000010000000000: n13731_o = 2'b00;
      15'b000001000000000: n13731_o = 2'b10;
      15'b000000100000000: n13731_o = 2'b01;
      15'b000000010000000: n13731_o = n13641_o;
      15'b000000001000000: n13731_o = 2'b10;
      15'b000000000100000: n13731_o = 2'b10;
      15'b000000000010000: n13731_o = 2'b10;
      15'b000000000001000: n13731_o = 2'b10;
      15'b000000000000100: n13731_o = 2'b00;
      15'b000000000000010: n13731_o = 2'b00;
      15'b000000000000001: n13731_o = n13588_o;
      default: n13731_o = 2'b00;
    endcase
  /* fpu.vhdl:784:21  */
  always @*
    case (n13717_o)
      15'b100000000000000: n13734_o = 1'b0;
      15'b010000000000000: n13734_o = 1'b0;
      15'b001000000000000: n13734_o = 1'b0;
      15'b000100000000000: n13734_o = 1'b0;
      15'b000010000000000: n13734_o = 1'b0;
      15'b000001000000000: n13734_o = 1'b0;
      15'b000000100000000: n13734_o = 1'b0;
      15'b000000010000000: n13734_o = 1'b0;
      15'b000000001000000: n13734_o = 1'b0;
      15'b000000000100000: n13734_o = 1'b0;
      15'b000000000010000: n13734_o = 1'b0;
      15'b000000000001000: n13734_o = 1'b0;
      15'b000000000000100: n13734_o = 1'b0;
      15'b000000000000010: n13734_o = 1'b0;
      15'b000000000000001: n13734_o = 1'b0;
      default: n13734_o = 1'b1;
    endcase
  assign n13735_o = {n13730_o, n13726_o};
  /* fpu.vhdl:783:17  */
  assign n13736_o = n13573_o ? n13718_o : n13151_o;
  assign n13737_o = n13465_o[5:3];
  assign n13738_o = r[702:700];
  /* fpu.vhdl:650:9  */
  assign n13739_o = n13152_o ? n13737_o : n13738_o;
  /* fpu.vhdl:783:17  */
  assign n13740_o = n13573_o ? n13722_o : n13739_o;
  assign n13741_o = n13465_o[11:10];
  assign n13742_o = r[708:707];
  /* fpu.vhdl:650:9  */
  assign n13743_o = n13152_o ? n13741_o : n13742_o;
  /* fpu.vhdl:783:17  */
  assign n13744_o = n13573_o ? n13735_o : n13743_o;
  /* fpu.vhdl:783:17  */
  assign n13745_o = n13573_o ? n13731_o : 2'b00;
  /* fpu.vhdl:783:17  */
  assign n13747_o = n13573_o ? n13734_o : 1'b0;
  /* fpu.vhdl:879:37  */
  assign n13749_o = r[156:152];
  /* fpu.vhdl:777:13  */
  assign n13751_o = n13567_o == 7'b0000000;
  /* fpu.vhdl:883:53  */
  assign n13753_o = r[48:17];
  /* insn_helpers.vhdl:141:23  */
  assign n13758_o = n13753_o[20:18];
  /* fpu.vhdl:883:22  */
  assign n13759_o = {28'b0, n13758_o};  //  uext
  /* fpu.vhdl:883:17  */
  assign n13760_o = {1'b0, n13759_o};  //  uext
  /* fpu.vhdl:885:26  */
  assign n13762_o = 32'b00000000000000000000000000000000 == n13760_o;
  /* fpu.vhdl:887:47  */
  assign n13763_o = r[158:155];
  /* fpu.vhdl:885:21  */
  assign n13765_o = n13762_o ? n13763_o : n13487_o;
  /* fpu.vhdl:885:21  */
  assign n13767_o = n13762_o ? 4'b0000 : 4'b1111;
  /* fpu.vhdl:885:26  */
  assign n13771_o = 32'b00000000000000000000000000000001 == n13760_o;
  /* fpu.vhdl:887:47  */
  assign n13772_o = r[154:151];
  /* fpu.vhdl:885:21  */
  assign n13774_o = n13771_o ? n13772_o : n13765_o;
  /* fpu.vhdl:885:21  */
  assign n13776_o = n13771_o ? 4'b0000 : 4'b1111;
  /* fpu.vhdl:885:26  */
  assign n13780_o = 32'b00000000000000000000000000000010 == n13760_o;
  /* fpu.vhdl:887:47  */
  assign n13781_o = r[150:147];
  /* fpu.vhdl:885:21  */
  assign n13783_o = n13780_o ? n13781_o : n13774_o;
  /* fpu.vhdl:885:21  */
  assign n13785_o = n13780_o ? 4'b0000 : 4'b1111;
  /* fpu.vhdl:885:26  */
  assign n13789_o = 32'b00000000000000000000000000000011 == n13760_o;
  /* fpu.vhdl:887:47  */
  assign n13790_o = r[146:143];
  /* fpu.vhdl:885:21  */
  assign n13792_o = n13789_o ? n13790_o : n13783_o;
  /* fpu.vhdl:885:21  */
  assign n13794_o = n13789_o ? 4'b0000 : 4'b1111;
  /* fpu.vhdl:885:26  */
  assign n13798_o = 32'b00000000000000000000000000000100 == n13760_o;
  /* fpu.vhdl:887:47  */
  assign n13799_o = r[142:139];
  /* fpu.vhdl:885:21  */
  assign n13801_o = n13798_o ? n13799_o : n13792_o;
  /* fpu.vhdl:885:21  */
  assign n13803_o = n13798_o ? 4'b0000 : 4'b1111;
  /* fpu.vhdl:885:26  */
  assign n13807_o = 32'b00000000000000000000000000000101 == n13760_o;
  /* fpu.vhdl:887:47  */
  assign n13808_o = r[138:135];
  /* fpu.vhdl:885:21  */
  assign n13810_o = n13807_o ? n13808_o : n13801_o;
  /* fpu.vhdl:885:21  */
  assign n13812_o = n13807_o ? 4'b0000 : 4'b1111;
  /* fpu.vhdl:885:26  */
  assign n13816_o = 32'b00000000000000000000000000000110 == n13760_o;
  /* fpu.vhdl:887:47  */
  assign n13817_o = r[134:131];
  /* fpu.vhdl:885:21  */
  assign n13819_o = n13816_o ? n13817_o : n13810_o;
  /* fpu.vhdl:885:21  */
  assign n13821_o = n13816_o ? 4'b0000 : 4'b1111;
  /* fpu.vhdl:885:26  */
  assign n13825_o = 32'b00000000000000000000000000000111 == n13760_o;
  /* fpu.vhdl:887:47  */
  assign n13826_o = r[130:127];
  /* fpu.vhdl:885:21  */
  assign n13828_o = n13825_o ? n13826_o : n13819_o;
  /* fpu.vhdl:885:21  */
  assign n13830_o = n13825_o ? 4'b0000 : 4'b1111;
  /* fpu.vhdl:891:30  */
  assign n13833_o = r[158:127];
  assign n13835_o = {n13767_o, n13776_o, n13785_o, n13794_o, n13803_o, n13812_o, n13821_o, n13830_o};
  /* fpu.vhdl:891:52  */
  assign n13836_o = n13835_o | 32'b01100000000001111111100011111111;
  /* fpu.vhdl:891:36  */
  assign n13837_o = n13833_o & n13836_o;
  /* fpu.vhdl:882:13  */
  assign n13841_o = n13567_o == 7'b0000001;
  /* fpu.vhdl:899:22  */
  assign n13845_o = r[238:159];
  /* fpu.vhdl:899:24  */
  assign n13846_o = n13845_o[1:0];
  /* fpu.vhdl:899:30  */
  assign n13848_o = n13846_o == 2'b10;
  /* fpu.vhdl:899:46  */
  assign n13849_o = r[318:239];
  /* fpu.vhdl:899:48  */
  assign n13850_o = n13849_o[1:0];
  /* fpu.vhdl:899:54  */
  assign n13852_o = n13850_o == 2'b00;
  /* fpu.vhdl:899:41  */
  assign n13853_o = n13848_o | n13852_o;
  /* fpu.vhdl:899:66  */
  assign n13854_o = r[318:239];
  /* fpu.vhdl:899:68  */
  assign n13855_o = n13854_o[1:0];
  /* fpu.vhdl:899:74  */
  assign n13857_o = n13855_o == 2'b10;
  /* fpu.vhdl:899:61  */
  assign n13858_o = n13853_o | n13857_o;
  /* fpu.vhdl:900:24  */
  assign n13859_o = r[318:239];
  /* fpu.vhdl:900:26  */
  assign n13860_o = n13859_o[1:0];
  /* fpu.vhdl:900:32  */
  assign n13862_o = n13860_o == 2'b01;
  /* fpu.vhdl:900:57  */
  assign n13863_o = r[308];
  /* fpu.vhdl:900:62  */
  assign n13864_o = ~n13863_o;
  /* fpu.vhdl:900:41  */
  assign n13865_o = n13862_o & n13864_o;
  /* fpu.vhdl:899:85  */
  assign n13866_o = n13858_o | n13865_o;
  assign n13868_o = n13844_o[2];
  /* fpu.vhdl:899:17  */
  assign n13869_o = n13866_o ? 1'b1 : n13868_o;
  assign n13870_o = n13844_o[3];
  /* fpu.vhdl:903:22  */
  assign n13872_o = r[238:159];
  /* fpu.vhdl:903:24  */
  assign n13873_o = n13872_o[1:0];
  /* fpu.vhdl:903:30  */
  assign n13875_o = n13873_o == 2'b11;
  /* fpu.vhdl:903:41  */
  assign n13876_o = r[238:159];
  /* fpu.vhdl:903:43  */
  assign n13877_o = n13876_o[1:0];
  /* fpu.vhdl:903:49  */
  assign n13879_o = n13877_o == 2'b10;
  /* fpu.vhdl:903:36  */
  assign n13880_o = n13875_o | n13879_o;
  /* fpu.vhdl:904:23  */
  assign n13881_o = r[318:239];
  /* fpu.vhdl:904:25  */
  assign n13882_o = n13881_o[1:0];
  /* fpu.vhdl:904:31  */
  assign n13884_o = n13882_o == 2'b11;
  /* fpu.vhdl:903:60  */
  assign n13885_o = n13880_o | n13884_o;
  /* fpu.vhdl:904:42  */
  assign n13886_o = r[318:239];
  /* fpu.vhdl:904:44  */
  assign n13887_o = n13886_o[1:0];
  /* fpu.vhdl:904:50  */
  assign n13889_o = n13887_o == 2'b00;
  /* fpu.vhdl:904:37  */
  assign n13890_o = n13885_o | n13889_o;
  /* fpu.vhdl:904:62  */
  assign n13891_o = r[318:239];
  /* fpu.vhdl:904:64  */
  assign n13892_o = n13891_o[1:0];
  /* fpu.vhdl:904:70  */
  assign n13894_o = n13892_o == 2'b10;
  /* fpu.vhdl:904:57  */
  assign n13895_o = n13890_o | n13894_o;
  /* fpu.vhdl:905:24  */
  assign n13896_o = r[238:159];
  /* fpu.vhdl:905:26  */
  assign n13897_o = n13896_o[1:0];
  /* fpu.vhdl:905:32  */
  assign n13899_o = n13897_o == 2'b01;
  /* fpu.vhdl:905:47  */
  assign n13900_o = r[238:159];
  /* fpu.vhdl:905:49  */
  assign n13901_o = n13900_o[15:3];
  /* fpu.vhdl:905:58  */
  assign n13903_o = $signed(n13901_o) <= $signed(13'b1110000110110);
  /* fpu.vhdl:905:41  */
  assign n13904_o = n13899_o & n13903_o;
  /* fpu.vhdl:904:81  */
  assign n13905_o = n13895_o | n13904_o;
  /* fpu.vhdl:903:17  */
  assign n13911_o = n13905_o ? 7'b0000000 : 7'b0101101;
  /* fpu.vhdl:903:17  */
  assign n13912_o = n13905_o ? 1'b1 : 1'b0;
  assign n13913_o = n13844_o[1];
  /* fpu.vhdl:903:17  */
  assign n13914_o = n13905_o ? 1'b1 : n13913_o;
  /* fpu.vhdl:903:17  */
  assign n13915_o = n13905_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:903:17  */
  assign n13916_o = n13905_o ? n13477_o : 2'b11;
  assign n13917_o = n13844_o[0];
  /* fpu.vhdl:895:13  */
  assign n13919_o = n13567_o == 7'b0001001;
  /* fpu.vhdl:918:22  */
  assign n13923_o = r[318:239];
  /* fpu.vhdl:918:24  */
  assign n13924_o = n13923_o[1:0];
  /* fpu.vhdl:918:30  */
  assign n13926_o = n13924_o == 2'b00;
  /* fpu.vhdl:918:42  */
  assign n13927_o = r[318:239];
  /* fpu.vhdl:918:44  */
  assign n13928_o = n13927_o[1:0];
  /* fpu.vhdl:918:50  */
  assign n13930_o = n13928_o == 2'b10;
  /* fpu.vhdl:918:37  */
  assign n13931_o = n13926_o | n13930_o;
  /* fpu.vhdl:919:24  */
  assign n13932_o = r[318:239];
  /* fpu.vhdl:919:26  */
  assign n13933_o = n13932_o[1:0];
  /* fpu.vhdl:919:32  */
  assign n13935_o = n13933_o == 2'b01;
  /* fpu.vhdl:919:57  */
  assign n13936_o = r[308];
  /* fpu.vhdl:919:62  */
  assign n13937_o = ~n13936_o;
  /* fpu.vhdl:919:41  */
  assign n13938_o = n13935_o & n13937_o;
  /* fpu.vhdl:918:61  */
  assign n13939_o = n13931_o | n13938_o;
  assign n13941_o = n13922_o[2];
  /* fpu.vhdl:918:17  */
  assign n13942_o = n13939_o ? 1'b1 : n13941_o;
  assign n13943_o = n13922_o[3];
  /* fpu.vhdl:922:22  */
  assign n13945_o = r[318:239];
  /* fpu.vhdl:922:24  */
  assign n13946_o = n13945_o[1:0];
  /* fpu.vhdl:922:30  */
  assign n13948_o = n13946_o == 2'b11;
  /* fpu.vhdl:922:41  */
  assign n13949_o = r[318:239];
  /* fpu.vhdl:922:43  */
  assign n13950_o = n13949_o[1:0];
  /* fpu.vhdl:922:49  */
  assign n13952_o = n13950_o == 2'b10;
  /* fpu.vhdl:922:36  */
  assign n13953_o = n13948_o | n13952_o;
  /* fpu.vhdl:922:65  */
  assign n13954_o = r[318:239];
  /* fpu.vhdl:922:67  */
  assign n13955_o = n13954_o[1:0];
  /* fpu.vhdl:922:73  */
  assign n13957_o = n13955_o == 2'b00;
  /* fpu.vhdl:922:60  */
  assign n13958_o = n13953_o | n13957_o;
  /* fpu.vhdl:923:26  */
  assign n13959_o = r[318:239];
  /* fpu.vhdl:923:28  */
  assign n13960_o = n13959_o[2];
  /* fpu.vhdl:923:21  */
  assign n13961_o = n13958_o | n13960_o;
  /* fpu.vhdl:923:48  */
  assign n13962_o = r[318:239];
  /* fpu.vhdl:923:50  */
  assign n13963_o = n13962_o[15:3];
  /* fpu.vhdl:923:59  */
  assign n13965_o = $signed(n13963_o) <= $signed(13'b1110000110110);
  /* fpu.vhdl:923:43  */
  assign n13966_o = n13961_o | n13965_o;
  assign n13968_o = n13922_o[1];
  /* fpu.vhdl:922:17  */
  assign n13969_o = n13966_o ? 1'b0 : n13968_o;
  assign n13970_o = n13922_o[0];
  /* fpu.vhdl:914:13  */
  assign n13972_o = n13567_o == 7'b0001010;
  /* fpu.vhdl:933:35  */
  assign n13975_o = r[318:239];
  /* fpu.vhdl:933:37  */
  assign n13976_o = n13975_o[15:3];
  /* fpu.vhdl:934:23  */
  assign n13977_o = r[238:159];
  /* fpu.vhdl:934:25  */
  assign n13978_o = n13977_o[1:0];
  /* fpu.vhdl:934:31  */
  assign n13980_o = n13978_o == 2'b11;
  /* fpu.vhdl:934:53  */
  assign n13981_o = r[228];
  /* fpu.vhdl:934:58  */
  assign n13982_o = ~n13981_o;
  /* fpu.vhdl:934:37  */
  assign n13983_o = n13980_o & n13982_o;
  /* fpu.vhdl:935:24  */
  assign n13984_o = r[318:239];
  /* fpu.vhdl:935:26  */
  assign n13985_o = n13984_o[1:0];
  /* fpu.vhdl:935:32  */
  assign n13987_o = n13985_o == 2'b11;
  /* fpu.vhdl:935:54  */
  assign n13988_o = r[308];
  /* fpu.vhdl:935:59  */
  assign n13989_o = ~n13988_o;
  /* fpu.vhdl:935:38  */
  assign n13990_o = n13987_o & n13989_o;
  /* fpu.vhdl:934:65  */
  assign n13991_o = n13983_o | n13990_o;
  /* fpu.vhdl:938:30  */
  assign n13993_o = r[23];
  /* fpu.vhdl:938:51  */
  assign n13994_o = r[134];
  /* fpu.vhdl:938:62  */
  assign n13995_o = ~n13994_o;
  /* fpu.vhdl:938:40  */
  assign n13996_o = n13993_o & n13995_o;
  assign n13998_o = r[146];
  /* fpu.vhdl:938:21  */
  assign n13999_o = n13996_o ? 1'b1 : n13998_o;
  /* fpu.vhdl:943:25  */
  assign n14001_o = r[238:159];
  /* fpu.vhdl:943:27  */
  assign n14002_o = n14001_o[1:0];
  /* fpu.vhdl:943:33  */
  assign n14004_o = n14002_o == 2'b11;
  /* fpu.vhdl:943:44  */
  assign n14005_o = r[318:239];
  /* fpu.vhdl:943:46  */
  assign n14006_o = n14005_o[1:0];
  /* fpu.vhdl:943:52  */
  assign n14008_o = n14006_o == 2'b11;
  /* fpu.vhdl:943:39  */
  assign n14009_o = n14004_o | n14008_o;
  /* fpu.vhdl:944:30  */
  assign n14010_o = r[23];
  assign n14012_o = r[146];
  /* fpu.vhdl:943:17  */
  assign n14013_o = n14155_o ? 1'b1 : n14012_o;
  /* fpu.vhdl:944:21  */
  assign n14016_o = n14010_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:950:25  */
  assign n14018_o = r[238:159];
  /* fpu.vhdl:950:27  */
  assign n14019_o = n14018_o[1:0];
  /* fpu.vhdl:950:33  */
  assign n14021_o = n14019_o == 2'b00;
  /* fpu.vhdl:950:46  */
  assign n14022_o = r[318:239];
  /* fpu.vhdl:950:48  */
  assign n14023_o = n14022_o[1:0];
  /* fpu.vhdl:950:54  */
  assign n14025_o = n14023_o == 2'b00;
  /* fpu.vhdl:950:40  */
  assign n14026_o = n14021_o & n14025_o;
  /* fpu.vhdl:952:25  */
  assign n14028_o = r[238:159];
  /* fpu.vhdl:952:27  */
  assign n14029_o = n14028_o[2];
  /* fpu.vhdl:952:41  */
  assign n14030_o = r[318:239];
  /* fpu.vhdl:952:43  */
  assign n14031_o = n14030_o[2];
  /* fpu.vhdl:952:36  */
  assign n14032_o = n14029_o != n14031_o;
  /* fpu.vhdl:953:38  */
  assign n14033_o = r[238:159];
  /* fpu.vhdl:953:40  */
  assign n14034_o = n14033_o[2];
  /* fpu.vhdl:953:53  */
  assign n14035_o = r[318:239];
  /* fpu.vhdl:953:55  */
  assign n14036_o = n14035_o[2];
  /* fpu.vhdl:953:49  */
  assign n14037_o = {n14034_o, n14036_o};
  /* fpu.vhdl:953:64  */
  assign n14039_o = {n14037_o, 2'b00};
  /* fpu.vhdl:954:25  */
  assign n14040_o = r[238:159];
  /* fpu.vhdl:954:27  */
  assign n14041_o = n14040_o[1:0];
  /* fpu.vhdl:954:33  */
  assign n14043_o = n14041_o == 2'b00;
  /* fpu.vhdl:956:42  */
  assign n14044_o = r[318:239];
  /* fpu.vhdl:956:44  */
  assign n14045_o = n14044_o[2];
  /* fpu.vhdl:956:36  */
  assign n14046_o = ~n14045_o;
  /* fpu.vhdl:956:57  */
  assign n14047_o = r[318:239];
  /* fpu.vhdl:956:59  */
  assign n14048_o = n14047_o[2];
  /* fpu.vhdl:956:53  */
  assign n14049_o = {n14046_o, n14048_o};
  /* fpu.vhdl:956:68  */
  assign n14051_o = {n14049_o, 2'b00};
  /* fpu.vhdl:957:25  */
  assign n14052_o = r[238:159];
  /* fpu.vhdl:957:27  */
  assign n14053_o = n14052_o[1:0];
  /* fpu.vhdl:957:33  */
  assign n14055_o = n14053_o == 2'b10;
  /* fpu.vhdl:958:26  */
  assign n14056_o = r[318:239];
  /* fpu.vhdl:958:28  */
  assign n14057_o = n14056_o[1:0];
  /* fpu.vhdl:958:34  */
  assign n14059_o = n14057_o == 2'b10;
  /* fpu.vhdl:961:42  */
  assign n14061_o = r[238:159];
  /* fpu.vhdl:961:44  */
  assign n14062_o = n14061_o[2];
  /* fpu.vhdl:961:61  */
  assign n14063_o = r[238:159];
  /* fpu.vhdl:961:63  */
  assign n14064_o = n14063_o[2];
  /* fpu.vhdl:961:55  */
  assign n14065_o = ~n14064_o;
  /* fpu.vhdl:961:53  */
  assign n14066_o = {n14062_o, n14065_o};
  /* fpu.vhdl:961:72  */
  assign n14068_o = {n14066_o, 2'b00};
  /* fpu.vhdl:958:21  */
  assign n14069_o = n14059_o ? 4'b0010 : n14068_o;
  /* fpu.vhdl:963:25  */
  assign n14070_o = r[318:239];
  /* fpu.vhdl:963:27  */
  assign n14071_o = n14070_o[1:0];
  /* fpu.vhdl:963:33  */
  assign n14073_o = n14071_o == 2'b00;
  /* fpu.vhdl:965:38  */
  assign n14074_o = r[238:159];
  /* fpu.vhdl:965:40  */
  assign n14075_o = n14074_o[2];
  /* fpu.vhdl:965:57  */
  assign n14076_o = r[238:159];
  /* fpu.vhdl:965:59  */
  assign n14077_o = n14076_o[2];
  /* fpu.vhdl:965:51  */
  assign n14078_o = ~n14077_o;
  /* fpu.vhdl:965:49  */
  assign n14079_o = {n14075_o, n14078_o};
  /* fpu.vhdl:965:68  */
  assign n14081_o = {n14079_o, 2'b00};
  /* fpu.vhdl:966:25  */
  assign n14082_o = r[318:239];
  /* fpu.vhdl:966:27  */
  assign n14083_o = n14082_o[1:0];
  /* fpu.vhdl:966:33  */
  assign n14085_o = n14083_o == 2'b10;
  /* fpu.vhdl:967:42  */
  assign n14086_o = r[318:239];
  /* fpu.vhdl:967:44  */
  assign n14087_o = n14086_o[2];
  /* fpu.vhdl:967:36  */
  assign n14088_o = ~n14087_o;
  /* fpu.vhdl:967:57  */
  assign n14089_o = r[318:239];
  /* fpu.vhdl:967:59  */
  assign n14090_o = n14089_o[2];
  /* fpu.vhdl:967:53  */
  assign n14091_o = {n14088_o, n14090_o};
  /* fpu.vhdl:967:68  */
  assign n14093_o = {n14091_o, 2'b00};
  /* fpu.vhdl:968:25  */
  assign n14094_o = r[704];
  /* fpu.vhdl:970:38  */
  assign n14095_o = r[238:159];
  /* fpu.vhdl:970:40  */
  assign n14096_o = n14095_o[2];
  /* fpu.vhdl:970:57  */
  assign n14097_o = r[238:159];
  /* fpu.vhdl:970:59  */
  assign n14098_o = n14097_o[2];
  /* fpu.vhdl:970:51  */
  assign n14099_o = ~n14098_o;
  /* fpu.vhdl:970:49  */
  assign n14100_o = {n14096_o, n14099_o};
  /* fpu.vhdl:970:68  */
  assign n14102_o = {n14100_o, 2'b00};
  /* fpu.vhdl:971:25  */
  assign n14103_o = r[238:159];
  /* fpu.vhdl:971:27  */
  assign n14104_o = n14103_o[15:3];
  /* fpu.vhdl:971:41  */
  assign n14105_o = r[318:239];
  /* fpu.vhdl:971:43  */
  assign n14106_o = n14105_o[15:3];
  /* fpu.vhdl:971:36  */
  assign n14107_o = n14104_o != n14106_o;
  /* fpu.vhdl:973:42  */
  assign n14108_o = r[238:159];
  /* fpu.vhdl:973:44  */
  assign n14109_o = n14108_o[2];
  /* fpu.vhdl:973:36  */
  assign n14110_o = ~n14109_o;
  /* fpu.vhdl:973:57  */
  assign n14111_o = r[238:159];
  /* fpu.vhdl:973:59  */
  assign n14112_o = n14111_o[2];
  /* fpu.vhdl:973:53  */
  assign n14113_o = {n14110_o, n14112_o};
  /* fpu.vhdl:973:68  */
  assign n14115_o = {n14113_o, 2'b00};
  /* fpu.vhdl:971:17  */
  assign n14120_o = n14107_o ? 7'b0000000 : 7'b0011100;
  /* fpu.vhdl:971:17  */
  assign n14121_o = n14107_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:971:17  */
  assign n14122_o = n14107_o ? n14115_o : 4'b0000;
  /* fpu.vhdl:971:17  */
  assign n14123_o = n14107_o ? 2'b00 : 2'b01;
  /* fpu.vhdl:968:17  */
  assign n14124_o = n14094_o ? 7'b0000000 : n14120_o;
  /* fpu.vhdl:968:17  */
  assign n14125_o = n14094_o ? 1'b1 : n14121_o;
  /* fpu.vhdl:968:17  */
  assign n14126_o = n14094_o ? n14102_o : n14122_o;
  /* fpu.vhdl:968:17  */
  assign n14127_o = n14094_o ? 2'b00 : n14123_o;
  /* fpu.vhdl:966:17  */
  assign n14128_o = n14085_o ? 7'b0000000 : n14124_o;
  /* fpu.vhdl:966:17  */
  assign n14129_o = n14085_o ? 1'b1 : n14125_o;
  /* fpu.vhdl:966:17  */
  assign n14130_o = n14085_o ? n14093_o : n14126_o;
  /* fpu.vhdl:966:17  */
  assign n14131_o = n14085_o ? 2'b00 : n14127_o;
  /* fpu.vhdl:963:17  */
  assign n14132_o = n14073_o ? 7'b0000000 : n14128_o;
  /* fpu.vhdl:963:17  */
  assign n14133_o = n14073_o ? 1'b1 : n14129_o;
  /* fpu.vhdl:963:17  */
  assign n14134_o = n14073_o ? n14081_o : n14130_o;
  /* fpu.vhdl:963:17  */
  assign n14135_o = n14073_o ? 2'b00 : n14131_o;
  /* fpu.vhdl:957:17  */
  assign n14136_o = n14055_o ? 7'b0000000 : n14132_o;
  /* fpu.vhdl:957:17  */
  assign n14137_o = n14055_o ? 1'b1 : n14133_o;
  /* fpu.vhdl:957:17  */
  assign n14138_o = n14055_o ? n14069_o : n14134_o;
  /* fpu.vhdl:957:17  */
  assign n14139_o = n14055_o ? 2'b00 : n14135_o;
  /* fpu.vhdl:954:17  */
  assign n14140_o = n14043_o ? 7'b0000000 : n14136_o;
  /* fpu.vhdl:954:17  */
  assign n14141_o = n14043_o ? 1'b1 : n14137_o;
  /* fpu.vhdl:954:17  */
  assign n14142_o = n14043_o ? n14051_o : n14138_o;
  /* fpu.vhdl:954:17  */
  assign n14143_o = n14043_o ? 2'b00 : n14139_o;
  /* fpu.vhdl:952:17  */
  assign n14144_o = n14032_o ? 7'b0000000 : n14140_o;
  /* fpu.vhdl:952:17  */
  assign n14145_o = n14032_o ? 1'b1 : n14141_o;
  /* fpu.vhdl:952:17  */
  assign n14146_o = n14032_o ? n14039_o : n14142_o;
  /* fpu.vhdl:952:17  */
  assign n14147_o = n14032_o ? 2'b00 : n14143_o;
  /* fpu.vhdl:950:17  */
  assign n14148_o = n14026_o ? 7'b0000000 : n14144_o;
  /* fpu.vhdl:950:17  */
  assign n14149_o = n14026_o ? 1'b1 : n14145_o;
  /* fpu.vhdl:950:17  */
  assign n14150_o = n14026_o ? 4'b0010 : n14146_o;
  /* fpu.vhdl:950:17  */
  assign n14151_o = n14026_o ? 2'b00 : n14147_o;
  /* fpu.vhdl:943:17  */
  assign n14152_o = n14009_o ? 7'b0000000 : n14148_o;
  /* fpu.vhdl:943:17  */
  assign n14153_o = n14009_o ? 1'b1 : n14149_o;
  /* fpu.vhdl:943:17  */
  assign n14155_o = n14009_o & n14010_o;
  /* fpu.vhdl:943:17  */
  assign n14156_o = n14009_o ? 4'b0001 : n14150_o;
  /* fpu.vhdl:943:17  */
  assign n14157_o = n14009_o ? 2'b00 : n14151_o;
  /* fpu.vhdl:943:17  */
  assign n14159_o = n14009_o ? n14016_o : 1'b0;
  /* fpu.vhdl:934:17  */
  assign n14160_o = n13991_o ? 7'b0000000 : n14152_o;
  /* fpu.vhdl:934:17  */
  assign n14161_o = n13991_o ? 1'b1 : n14153_o;
  /* fpu.vhdl:934:17  */
  assign n14162_o = n13991_o ? n13999_o : n14013_o;
  assign n14163_o = r[151];
  /* fpu.vhdl:934:17  */
  assign n14164_o = n13991_o ? 1'b1 : n14163_o;
  /* fpu.vhdl:934:17  */
  assign n14165_o = n13991_o ? 4'b0001 : n14156_o;
  /* fpu.vhdl:934:17  */
  assign n14166_o = n13991_o ? 2'b00 : n14157_o;
  /* fpu.vhdl:934:17  */
  assign n14168_o = n13991_o ? 1'b1 : n14159_o;
  assign n14169_o = r[145:127];
  assign n14170_o = r[150:147];
  assign n14171_o = r[158:152];
  assign n14172_o = r[650:399];
  assign n14173_o = {n13479_o, n13564_o, n14166_o, n13477_o, n13562_o, 1'b0, n13475_o, 1'b0, n13558_o, n13473_o, n14165_o, n13471_o, 1'b0, 13'b0000000000000, n13976_o, n14172_o, n13469_o, n14171_o, n14164_o, n14170_o, n14162_o, n14169_o, n13467_o, n13556_o, n14161_o, 1'b0, n14160_o};
  /* fpu.vhdl:981:56  */
  assign n14174_o = n14173_o[682:679];
  /* fpu.vhdl:927:13  */
  assign n14176_o = n13567_o == 7'b0001000;
  /* fpu.vhdl:985:52  */
  assign n14178_o = r[48:17];
  /* insn_helpers.vhdl:161:23  */
  assign n14183_o = n14178_o[25:21];
  /* fpu.vhdl:985:22  */
  assign n14184_o = {26'b0, n14183_o};  //  uext
  /* fpu.vhdl:985:17  */
  assign n14185_o = {1'b0, n14184_o};  //  uext
  /* fpu.vhdl:987:26  */
  assign n14187_o = 32'b00000000000000000000000000000000 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14188_o = r[23];
  assign n14189_o = r[158];
  /* fpu.vhdl:987:21  */
  assign n14190_o = n14187_o ? n14188_o : n14189_o;
  /* fpu.vhdl:987:26  */
  assign n14192_o = 32'b00000000000000000000000000000001 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14193_o = r[23];
  assign n14194_o = r[157];
  /* fpu.vhdl:987:21  */
  assign n14195_o = n14192_o ? n14193_o : n14194_o;
  /* fpu.vhdl:987:26  */
  assign n14197_o = 32'b00000000000000000000000000000010 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14198_o = r[23];
  assign n14199_o = r[156];
  /* fpu.vhdl:987:21  */
  assign n14200_o = n14197_o ? n14198_o : n14199_o;
  /* fpu.vhdl:987:26  */
  assign n14202_o = 32'b00000000000000000000000000000011 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14203_o = r[23];
  assign n14204_o = r[155];
  /* fpu.vhdl:987:21  */
  assign n14205_o = n14202_o ? n14203_o : n14204_o;
  /* fpu.vhdl:987:26  */
  assign n14207_o = 32'b00000000000000000000000000000100 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14208_o = r[23];
  assign n14209_o = r[154];
  /* fpu.vhdl:987:21  */
  assign n14210_o = n14207_o ? n14208_o : n14209_o;
  /* fpu.vhdl:987:26  */
  assign n14212_o = 32'b00000000000000000000000000000101 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14213_o = r[23];
  assign n14214_o = r[153];
  /* fpu.vhdl:987:21  */
  assign n14215_o = n14212_o ? n14213_o : n14214_o;
  /* fpu.vhdl:987:26  */
  assign n14217_o = 32'b00000000000000000000000000000110 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14218_o = r[23];
  assign n14219_o = r[152];
  /* fpu.vhdl:987:21  */
  assign n14220_o = n14217_o ? n14218_o : n14219_o;
  /* fpu.vhdl:987:26  */
  assign n14222_o = 32'b00000000000000000000000000000111 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14223_o = r[23];
  assign n14224_o = r[151];
  /* fpu.vhdl:987:21  */
  assign n14225_o = n14222_o ? n14223_o : n14224_o;
  /* fpu.vhdl:987:26  */
  assign n14227_o = 32'b00000000000000000000000000001000 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14228_o = r[23];
  assign n14229_o = r[150];
  /* fpu.vhdl:987:21  */
  assign n14230_o = n14227_o ? n14228_o : n14229_o;
  /* fpu.vhdl:987:26  */
  assign n14232_o = 32'b00000000000000000000000000001001 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14233_o = r[23];
  assign n14234_o = r[149];
  /* fpu.vhdl:987:21  */
  assign n14235_o = n14232_o ? n14233_o : n14234_o;
  /* fpu.vhdl:987:26  */
  assign n14237_o = 32'b00000000000000000000000000001010 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14238_o = r[23];
  assign n14239_o = r[148];
  /* fpu.vhdl:987:21  */
  assign n14240_o = n14237_o ? n14238_o : n14239_o;
  /* fpu.vhdl:987:26  */
  assign n14242_o = 32'b00000000000000000000000000001011 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14243_o = r[23];
  assign n14244_o = r[147];
  /* fpu.vhdl:987:21  */
  assign n14245_o = n14242_o ? n14243_o : n14244_o;
  /* fpu.vhdl:987:26  */
  assign n14247_o = 32'b00000000000000000000000000001100 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14248_o = r[23];
  assign n14249_o = r[146];
  /* fpu.vhdl:987:21  */
  assign n14250_o = n14247_o ? n14248_o : n14249_o;
  /* fpu.vhdl:987:26  */
  assign n14252_o = 32'b00000000000000000000000000001101 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14253_o = r[23];
  assign n14254_o = r[145];
  /* fpu.vhdl:987:21  */
  assign n14255_o = n14252_o ? n14253_o : n14254_o;
  /* fpu.vhdl:987:26  */
  assign n14257_o = 32'b00000000000000000000000000001110 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14258_o = r[23];
  assign n14259_o = r[144];
  /* fpu.vhdl:987:21  */
  assign n14260_o = n14257_o ? n14258_o : n14259_o;
  /* fpu.vhdl:987:26  */
  assign n14262_o = 32'b00000000000000000000000000001111 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14263_o = r[23];
  assign n14264_o = r[143];
  /* fpu.vhdl:987:21  */
  assign n14265_o = n14262_o ? n14263_o : n14264_o;
  /* fpu.vhdl:987:26  */
  assign n14267_o = 32'b00000000000000000000000000010000 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14268_o = r[23];
  assign n14269_o = r[142];
  /* fpu.vhdl:987:21  */
  assign n14270_o = n14267_o ? n14268_o : n14269_o;
  /* fpu.vhdl:987:26  */
  assign n14272_o = 32'b00000000000000000000000000010001 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14273_o = r[23];
  assign n14274_o = r[141];
  /* fpu.vhdl:987:21  */
  assign n14275_o = n14272_o ? n14273_o : n14274_o;
  /* fpu.vhdl:987:26  */
  assign n14277_o = 32'b00000000000000000000000000010010 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14278_o = r[23];
  assign n14279_o = r[140];
  /* fpu.vhdl:987:21  */
  assign n14280_o = n14277_o ? n14278_o : n14279_o;
  /* fpu.vhdl:987:26  */
  assign n14282_o = 32'b00000000000000000000000000010011 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14283_o = r[23];
  assign n14284_o = r[139];
  /* fpu.vhdl:987:21  */
  assign n14285_o = n14282_o ? n14283_o : n14284_o;
  /* fpu.vhdl:987:26  */
  assign n14287_o = 32'b00000000000000000000000000010100 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14288_o = r[23];
  assign n14289_o = r[138];
  /* fpu.vhdl:987:21  */
  assign n14290_o = n14287_o ? n14288_o : n14289_o;
  /* fpu.vhdl:987:26  */
  assign n14292_o = 32'b00000000000000000000000000010101 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14293_o = r[23];
  assign n14294_o = r[137];
  /* fpu.vhdl:987:21  */
  assign n14295_o = n14292_o ? n14293_o : n14294_o;
  /* fpu.vhdl:987:26  */
  assign n14297_o = 32'b00000000000000000000000000010110 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14298_o = r[23];
  assign n14299_o = r[136];
  /* fpu.vhdl:987:21  */
  assign n14300_o = n14297_o ? n14298_o : n14299_o;
  /* fpu.vhdl:987:26  */
  assign n14302_o = 32'b00000000000000000000000000010111 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14303_o = r[23];
  assign n14304_o = r[135];
  /* fpu.vhdl:987:21  */
  assign n14305_o = n14302_o ? n14303_o : n14304_o;
  /* fpu.vhdl:987:26  */
  assign n14307_o = 32'b00000000000000000000000000011000 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14308_o = r[23];
  assign n14309_o = r[134];
  /* fpu.vhdl:987:21  */
  assign n14310_o = n14307_o ? n14308_o : n14309_o;
  /* fpu.vhdl:987:26  */
  assign n14312_o = 32'b00000000000000000000000000011001 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14313_o = r[23];
  assign n14314_o = r[133];
  /* fpu.vhdl:987:21  */
  assign n14315_o = n14312_o ? n14313_o : n14314_o;
  /* fpu.vhdl:987:26  */
  assign n14317_o = 32'b00000000000000000000000000011010 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14318_o = r[23];
  assign n14319_o = r[132];
  /* fpu.vhdl:987:21  */
  assign n14320_o = n14317_o ? n14318_o : n14319_o;
  /* fpu.vhdl:987:26  */
  assign n14322_o = 32'b00000000000000000000000000011011 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14323_o = r[23];
  assign n14324_o = r[131];
  /* fpu.vhdl:987:21  */
  assign n14325_o = n14322_o ? n14323_o : n14324_o;
  /* fpu.vhdl:987:26  */
  assign n14327_o = 32'b00000000000000000000000000011100 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14328_o = r[23];
  assign n14329_o = r[130];
  /* fpu.vhdl:987:21  */
  assign n14330_o = n14327_o ? n14328_o : n14329_o;
  /* fpu.vhdl:987:26  */
  assign n14332_o = 32'b00000000000000000000000000011101 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14333_o = r[23];
  assign n14334_o = r[129];
  /* fpu.vhdl:987:21  */
  assign n14335_o = n14332_o ? n14333_o : n14334_o;
  /* fpu.vhdl:987:26  */
  assign n14337_o = 32'b00000000000000000000000000011110 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14338_o = r[23];
  assign n14339_o = r[128];
  /* fpu.vhdl:987:21  */
  assign n14340_o = n14337_o ? n14338_o : n14339_o;
  /* fpu.vhdl:987:26  */
  assign n14342_o = 32'b00000000000000000000000000011111 == n14185_o;
  /* fpu.vhdl:988:50  */
  assign n14343_o = r[23];
  assign n14344_o = r[127];
  /* fpu.vhdl:987:21  */
  assign n14345_o = n14342_o ? n14343_o : n14344_o;
  /* fpu.vhdl:983:13  */
  assign n14349_o = n13567_o == 7'b0000010;
  /* fpu.vhdl:996:52  */
  assign n14351_o = r[48:17];
  /* insn_helpers.vhdl:136:23  */
  assign n14356_o = n14351_o[25:23];
  /* fpu.vhdl:996:22  */
  assign n14357_o = {28'b0, n14356_o};  //  uext
  /* fpu.vhdl:996:17  */
  assign n14358_o = {1'b0, n14357_o};  //  uext
  /* fpu.vhdl:997:26  */
  assign n14359_o = r[33];
  /* fpu.vhdl:997:31  */
  assign n14360_o = ~n14359_o;
  /* fpu.vhdl:999:30  */
  assign n14362_o = 32'b00000000000000000000000000000000 == n14358_o;
  /* fpu.vhdl:1001:65  */
  assign n14364_o = r[48:17];
  /* insn_helpers.vhdl:251:23  */
  assign n14369_o = n14364_o[15:12];
  assign n14370_o = r[158:155];
  /* fpu.vhdl:999:25  */
  assign n14371_o = n14362_o ? n14369_o : n14370_o;
  /* fpu.vhdl:999:30  */
  assign n14375_o = 32'b00000000000000000000000000000001 == n14358_o;
  /* fpu.vhdl:1001:65  */
  assign n14377_o = r[48:17];
  /* insn_helpers.vhdl:251:23  */
  assign n14382_o = n14377_o[15:12];
  assign n14383_o = r[154:151];
  /* fpu.vhdl:999:25  */
  assign n14384_o = n14375_o ? n14382_o : n14383_o;
  /* fpu.vhdl:999:30  */
  assign n14388_o = 32'b00000000000000000000000000000010 == n14358_o;
  /* fpu.vhdl:1001:65  */
  assign n14390_o = r[48:17];
  /* insn_helpers.vhdl:251:23  */
  assign n14395_o = n14390_o[15:12];
  assign n14396_o = r[150:147];
  /* fpu.vhdl:999:25  */
  assign n14397_o = n14388_o ? n14395_o : n14396_o;
  /* fpu.vhdl:999:30  */
  assign n14401_o = 32'b00000000000000000000000000000011 == n14358_o;
  /* fpu.vhdl:1001:65  */
  assign n14403_o = r[48:17];
  /* insn_helpers.vhdl:251:23  */
  assign n14408_o = n14403_o[15:12];
  assign n14409_o = r[146:143];
  /* fpu.vhdl:999:25  */
  assign n14410_o = n14401_o ? n14408_o : n14409_o;
  /* fpu.vhdl:999:30  */
  assign n14414_o = 32'b00000000000000000000000000000100 == n14358_o;
  /* fpu.vhdl:1001:65  */
  assign n14416_o = r[48:17];
  /* insn_helpers.vhdl:251:23  */
  assign n14421_o = n14416_o[15:12];
  assign n14422_o = r[142:139];
  /* fpu.vhdl:999:25  */
  assign n14423_o = n14414_o ? n14421_o : n14422_o;
  /* fpu.vhdl:999:30  */
  assign n14427_o = 32'b00000000000000000000000000000101 == n14358_o;
  /* fpu.vhdl:1001:65  */
  assign n14429_o = r[48:17];
  /* insn_helpers.vhdl:251:23  */
  assign n14434_o = n14429_o[15:12];
  assign n14435_o = r[138:135];
  /* fpu.vhdl:999:25  */
  assign n14436_o = n14427_o ? n14434_o : n14435_o;
  /* fpu.vhdl:999:30  */
  assign n14440_o = 32'b00000000000000000000000000000110 == n14358_o;
  /* fpu.vhdl:1001:65  */
  assign n14442_o = r[48:17];
  /* insn_helpers.vhdl:251:23  */
  assign n14447_o = n14442_o[15:12];
  assign n14448_o = r[134:131];
  /* fpu.vhdl:999:25  */
  assign n14449_o = n14440_o ? n14447_o : n14448_o;
  /* fpu.vhdl:999:30  */
  assign n14453_o = 32'b00000000000000000000000000000111 == n14358_o;
  /* fpu.vhdl:1001:65  */
  assign n14455_o = r[48:17];
  /* insn_helpers.vhdl:251:23  */
  assign n14460_o = n14455_o[15:12];
  assign n14461_o = r[130:127];
  /* fpu.vhdl:999:25  */
  assign n14462_o = n14453_o ? n14460_o : n14461_o;
  assign n14465_o = {n14371_o, n14384_o, n14397_o, n14410_o, n14423_o, n14436_o, n14449_o, n14462_o};
  /* fpu.vhdl:997:17  */
  assign n14466_o = n14360_o ? n14465_o : n13483_o;
  /* fpu.vhdl:994:13  */
  assign n14471_o = n13567_o == 7'b0000011;
  /* fpu.vhdl:1011:42  */
  assign n14472_o = r[25];
  /* fpu.vhdl:1011:34  */
  assign n14474_o = {2'b01, n14472_o};
  /* fpu.vhdl:1011:46  */
  assign n14476_o = {n14474_o, 1'b0};
  /* fpu.vhdl:1008:13  */
  assign n14482_o = n13567_o == 7'b0000111;
  /* fpu.vhdl:1021:28  */
  assign n14485_o = r[37:33];
  /* fpu.vhdl:1022:21  */
  assign n14487_o = n14485_o == 5'b00000;
  /* fpu.vhdl:1024:21  */
  assign n14490_o = n14485_o == 5'b00001;
  /* fpu.vhdl:1027:21  */
  assign n14492_o = n14485_o == 5'b10100;
  /* fpu.vhdl:1027:34  */
  assign n14494_o = n14485_o == 5'b10101;
  /* fpu.vhdl:1027:34  */
  assign n14495_o = n14492_o | n14494_o;
  /* fpu.vhdl:1034:41  */
  assign n14496_o = r[256:255];
  /* fpu.vhdl:1030:21  */
  assign n14498_o = n14485_o == 5'b10110;
  /* fpu.vhdl:1038:70  */
  assign n14499_o = r[29:28];
  /* fpu.vhdl:1035:21  */
  assign n14501_o = n14485_o == 5'b10111;
  /* fpu.vhdl:1039:21  */
  assign n14503_o = n14485_o == 5'b11000;
  assign n14504_o = {n14503_o, n14501_o, n14498_o, n14495_o, n14490_o, n14487_o};
  assign n14505_o = r[128:127];
  /* fpu.vhdl:1021:17  */
  always @*
    case (n14504_o)
      6'b100000: n14506_o = n14505_o;
      6'b010000: n14506_o = n14499_o;
      6'b001000: n14506_o = n14496_o;
      6'b000100: n14506_o = n14505_o;
      6'b000010: n14506_o = n14505_o;
      6'b000001: n14506_o = n14505_o;
      default: n14506_o = n14505_o;
    endcase
  assign n14507_o = r[134:130];
  /* fpu.vhdl:1021:17  */
  always @*
    case (n14504_o)
      6'b100000: n14508_o = n14507_o;
      6'b010000: n14508_o = n14507_o;
      6'b001000: n14508_o = n14507_o;
      6'b000100: n14508_o = n14507_o;
      6'b000010: n14508_o = 5'b00000;
      6'b000001: n14508_o = n14507_o;
      default: n14508_o = n14507_o;
    endcase
  /* fpu.vhdl:1021:17  */
  always @*
    case (n14504_o)
      6'b100000: n14514_o = 32'b00000000000001111111000011111111;
      6'b010000: n14514_o = 32'b00000000000000000000000011111111;
      6'b001000: n14514_o = 32'b00000000000000000000000011111111;
      6'b000100: n14514_o = 32'b00000000000000000000000011111111;
      6'b000010: n14514_o = 32'b11111111111111111111111111111111;
      6'b000001: n14514_o = 32'b11111111111111111111111111111111;
      default: n14514_o = 32'b11111111111111111111111111111111;
    endcase
  /* fpu.vhdl:1021:17  */
  always @*
    case (n14504_o)
      6'b100000: n14517_o = 1'b0;
      6'b010000: n14517_o = 1'b0;
      6'b001000: n14517_o = 1'b0;
      6'b000100: n14517_o = 1'b0;
      6'b000010: n14517_o = 1'b0;
      6'b000001: n14517_o = 1'b0;
      default: n14517_o = 1'b1;
    endcase
  /* fpu.vhdl:1017:13  */
  assign n14521_o = n13567_o == 7'b0000100;
  /* fpu.vhdl:1049:26  */
  assign n14522_o = r[42];
  /* fpu.vhdl:1051:29  */
  assign n14523_o = r[33];
  /* fpu.vhdl:1054:34  */
  assign n14524_o = r[41:34];
  /* fpu.vhdl:1051:17  */
  assign n14526_o = n14523_o ? 8'b00000000 : n14524_o;
  /* fpu.vhdl:1049:17  */
  assign n14528_o = n14522_o ? 8'b11111111 : n14526_o;
  /* fpu.vhdl:1058:27  */
  assign n14529_o = n14528_o[0];
  /* fpu.vhdl:1059:64  */
  assign n14530_o = r[258:255];
  assign n14531_o = r[130:127];
  /* fpu.vhdl:1058:21  */
  assign n14532_o = n14529_o ? n14530_o : n14531_o;
  /* fpu.vhdl:1058:27  */
  assign n14533_o = n14528_o[1];
  /* fpu.vhdl:1059:64  */
  assign n14534_o = r[262:259];
  assign n14535_o = r[134:131];
  /* fpu.vhdl:1058:21  */
  assign n14536_o = n14533_o ? n14534_o : n14535_o;
  /* fpu.vhdl:1058:27  */
  assign n14537_o = n14528_o[2];
  /* fpu.vhdl:1059:64  */
  assign n14538_o = r[266:263];
  assign n14539_o = r[138:135];
  /* fpu.vhdl:1058:21  */
  assign n14540_o = n14537_o ? n14538_o : n14539_o;
  /* fpu.vhdl:1058:27  */
  assign n14541_o = n14528_o[3];
  /* fpu.vhdl:1059:64  */
  assign n14542_o = r[270:267];
  assign n14543_o = r[142:139];
  /* fpu.vhdl:1058:21  */
  assign n14544_o = n14541_o ? n14542_o : n14543_o;
  /* fpu.vhdl:1058:27  */
  assign n14545_o = n14528_o[4];
  /* fpu.vhdl:1059:64  */
  assign n14546_o = r[274:271];
  assign n14547_o = r[146:143];
  /* fpu.vhdl:1058:21  */
  assign n14548_o = n14545_o ? n14546_o : n14547_o;
  /* fpu.vhdl:1058:27  */
  assign n14549_o = n14528_o[5];
  /* fpu.vhdl:1059:64  */
  assign n14550_o = r[278:275];
  assign n14551_o = r[150:147];
  /* fpu.vhdl:1058:21  */
  assign n14552_o = n14549_o ? n14550_o : n14551_o;
  /* fpu.vhdl:1058:27  */
  assign n14553_o = n14528_o[6];
  /* fpu.vhdl:1059:64  */
  assign n14554_o = r[282:279];
  assign n14555_o = r[154:151];
  /* fpu.vhdl:1058:21  */
  assign n14556_o = n14553_o ? n14554_o : n14555_o;
  /* fpu.vhdl:1058:27  */
  assign n14557_o = n14528_o[7];
  /* fpu.vhdl:1059:64  */
  assign n14558_o = r[286:283];
  assign n14559_o = r[158:155];
  /* fpu.vhdl:1058:21  */
  assign n14560_o = n14557_o ? n14558_o : n14559_o;
  /* fpu.vhdl:1048:13  */
  assign n14564_o = n13567_o == 7'b0000101;
  /* fpu.vhdl:1067:37  */
  assign n14565_o = r[318:239];
  /* fpu.vhdl:1067:39  */
  assign n14566_o = n14565_o[1:0];
  /* fpu.vhdl:1068:35  */
  assign n14567_o = r[318:239];
  /* fpu.vhdl:1068:37  */
  assign n14568_o = n14567_o[15:3];
  /* fpu.vhdl:1070:26  */
  assign n14570_o = r[26];
  /* fpu.vhdl:1072:29  */
  assign n14572_o = r[25];
  /* fpu.vhdl:1074:29  */
  assign n14574_o = r[24];
  /* fpu.vhdl:1075:40  */
  assign n14575_o = r[318:239];
  /* fpu.vhdl:1075:42  */
  assign n14576_o = n14575_o[2];
  /* fpu.vhdl:1076:29  */
  assign n14577_o = r[23];
  /* fpu.vhdl:1077:44  */
  assign n14578_o = r[318:239];
  /* fpu.vhdl:1077:46  */
  assign n14579_o = n14578_o[2];
  /* fpu.vhdl:1077:38  */
  assign n14580_o = ~n14579_o;
  /* fpu.vhdl:1079:40  */
  assign n14581_o = r[238:159];
  /* fpu.vhdl:1079:42  */
  assign n14582_o = n14581_o[2];
  /* fpu.vhdl:1076:17  */
  assign n14583_o = n14577_o ? n14580_o : n14582_o;
  /* fpu.vhdl:1074:17  */
  assign n14584_o = n14574_o ? n14576_o : n14583_o;
  /* fpu.vhdl:1072:17  */
  assign n14585_o = n14572_o ? 1'b1 : n14584_o;
  /* fpu.vhdl:1070:17  */
  assign n14586_o = n14570_o ? 1'b0 : n14585_o;
  /* fpu.vhdl:1065:13  */
  assign n14591_o = n13567_o == 7'b0000110;
  /* fpu.vhdl:1087:37  */
  assign n14592_o = r[318:239];
  /* fpu.vhdl:1087:39  */
  assign n14593_o = n14592_o[1:0];
  /* fpu.vhdl:1088:36  */
  assign n14594_o = r[318:239];
  /* fpu.vhdl:1088:38  */
  assign n14595_o = n14594_o[2];
  /* fpu.vhdl:1089:35  */
  assign n14596_o = r[318:239];
  /* fpu.vhdl:1089:37  */
  assign n14597_o = n14596_o[15:3];
  /* fpu.vhdl:1092:22  */
  assign n14600_o = r[318:239];
  /* fpu.vhdl:1092:24  */
  assign n14601_o = n14600_o[1:0];
  /* fpu.vhdl:1092:30  */
  assign n14603_o = n14601_o == 2'b11;
  /* fpu.vhdl:1092:52  */
  assign n14604_o = r[308];
  /* fpu.vhdl:1092:57  */
  assign n14605_o = ~n14604_o;
  /* fpu.vhdl:1092:36  */
  assign n14606_o = n14603_o & n14605_o;
  assign n14608_o = r[151];
  /* fpu.vhdl:1092:17  */
  assign n14609_o = n14606_o ? 1'b1 : n14608_o;
  /* fpu.vhdl:1092:17  */
  assign n14612_o = n14606_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1097:22  */
  assign n14613_o = r[318:239];
  /* fpu.vhdl:1097:24  */
  assign n14614_o = n14613_o[1:0];
  /* fpu.vhdl:1097:30  */
  assign n14616_o = n14614_o == 2'b01;
  /* fpu.vhdl:1098:26  */
  assign n14617_o = r[318:239];
  /* fpu.vhdl:1098:28  */
  assign n14618_o = n14617_o[15:3];
  /* fpu.vhdl:1098:37  */
  assign n14620_o = $signed(n14618_o) >= $signed(13'b0000000110100);
  /* fpu.vhdl:1102:38  */
  assign n14621_o = r[318:239];
  /* fpu.vhdl:1102:40  */
  assign n14622_o = n14621_o[15:3];
  /* fpu.vhdl:1102:49  */
  assign n14624_o = n14622_o - 13'b0000000110100;
  /* fpu.vhdl:1104:53  */
  assign n14626_o = r[24:23];
  /* fpu.vhdl:1104:45  */
  assign n14628_o = {1'b1, n14626_o};
  /* fpu.vhdl:1098:21  */
  assign n14629_o = n14620_o ? n13151_o : 7'b0010111;
  /* fpu.vhdl:1098:21  */
  assign n14630_o = n14620_o ? 13'b0000000000000 : n14624_o;
  assign n14631_o = n13465_o[5:3];
  assign n14632_o = r[702:700];
  /* fpu.vhdl:650:9  */
  assign n14633_o = n13152_o ? n14631_o : n14632_o;
  /* fpu.vhdl:1098:21  */
  assign n14634_o = n14620_o ? n14633_o : n14628_o;
  /* fpu.vhdl:1098:21  */
  assign n14637_o = n14620_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1097:17  */
  assign n14638_o = n14616_o ? n14629_o : n13151_o;
  /* fpu.vhdl:1097:17  */
  assign n14639_o = n14616_o ? n14630_o : 13'b0000000000000;
  assign n14640_o = n13465_o[5:3];
  assign n14641_o = r[702:700];
  /* fpu.vhdl:650:9  */
  assign n14642_o = n13152_o ? n14640_o : n14641_o;
  /* fpu.vhdl:1097:17  */
  assign n14643_o = n14616_o ? n14634_o : n14642_o;
  /* fpu.vhdl:1097:17  */
  assign n14645_o = n14616_o ? n14637_o : 1'b1;
  /* fpu.vhdl:1085:13  */
  assign n14647_o = n13567_o == 7'b0001110;
  /* fpu.vhdl:1112:37  */
  assign n14648_o = r[318:239];
  /* fpu.vhdl:1112:39  */
  assign n14649_o = n14648_o[1:0];
  /* fpu.vhdl:1113:36  */
  assign n14650_o = r[318:239];
  /* fpu.vhdl:1113:38  */
  assign n14651_o = n14650_o[2];
  /* fpu.vhdl:1114:35  */
  assign n14652_o = r[318:239];
  /* fpu.vhdl:1114:37  */
  assign n14653_o = n14652_o[15:3];
  /* fpu.vhdl:1117:22  */
  assign n14656_o = r[318:239];
  /* fpu.vhdl:1117:24  */
  assign n14657_o = n14656_o[1:0];
  /* fpu.vhdl:1117:30  */
  assign n14659_o = n14657_o == 2'b11;
  /* fpu.vhdl:1117:52  */
  assign n14660_o = r[308];
  /* fpu.vhdl:1117:57  */
  assign n14661_o = ~n14660_o;
  /* fpu.vhdl:1117:36  */
  assign n14662_o = n14659_o & n14661_o;
  assign n14664_o = r[151];
  /* fpu.vhdl:1117:17  */
  assign n14665_o = n14662_o ? 1'b1 : n14664_o;
  /* fpu.vhdl:1117:17  */
  assign n14668_o = n14662_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1123:22  */
  assign n14669_o = r[318:239];
  /* fpu.vhdl:1123:24  */
  assign n14670_o = n14669_o[1:0];
  /* fpu.vhdl:1123:30  */
  assign n14672_o = n14670_o == 2'b01;
  /* fpu.vhdl:1124:26  */
  assign n14673_o = r[318:239];
  /* fpu.vhdl:1124:28  */
  assign n14674_o = n14673_o[15:3];
  /* fpu.vhdl:1124:37  */
  assign n14676_o = $signed(n14674_o) < $signed(13'b1111110000010);
  /* fpu.vhdl:1125:38  */
  assign n14677_o = r[318:239];
  /* fpu.vhdl:1125:40  */
  assign n14678_o = n14677_o[15:3];
  /* fpu.vhdl:1125:49  */
  assign n14680_o = n14678_o - 13'b1111110000010;
  /* fpu.vhdl:1127:29  */
  assign n14682_o = r[318:239];
  /* fpu.vhdl:1127:31  */
  assign n14683_o = n14682_o[15:3];
  /* fpu.vhdl:1127:40  */
  assign n14685_o = $signed(n14683_o) > $signed(13'b0000001111111);
  /* fpu.vhdl:1127:21  */
  assign n14688_o = n14685_o ? 7'b1000011 : 7'b1000100;
  /* fpu.vhdl:1124:21  */
  assign n14689_o = n14676_o ? 7'b1000010 : n14688_o;
  /* fpu.vhdl:1123:17  */
  assign n14690_o = n14692_o ? n14680_o : 13'b0000000000000;
  /* fpu.vhdl:1123:17  */
  assign n14691_o = n14672_o ? n14689_o : n13151_o;
  /* fpu.vhdl:1123:17  */
  assign n14692_o = n14672_o & n14676_o;
  /* fpu.vhdl:1123:17  */
  assign n14695_o = n14672_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:1110:13  */
  assign n14697_o = n13567_o == 7'b0001101;
  /* fpu.vhdl:1141:37  */
  assign n14698_o = r[318:239];
  /* fpu.vhdl:1141:39  */
  assign n14699_o = n14698_o[1:0];
  /* fpu.vhdl:1142:36  */
  assign n14700_o = r[318:239];
  /* fpu.vhdl:1142:38  */
  assign n14701_o = n14700_o[2];
  /* fpu.vhdl:1143:35  */
  assign n14702_o = r[318:239];
  /* fpu.vhdl:1143:37  */
  assign n14703_o = n14702_o[15:3];
  /* fpu.vhdl:1146:22  */
  assign n14706_o = r[318:239];
  /* fpu.vhdl:1146:24  */
  assign n14707_o = n14706_o[1:0];
  /* fpu.vhdl:1146:30  */
  assign n14709_o = n14707_o == 2'b11;
  /* fpu.vhdl:1146:52  */
  assign n14710_o = r[308];
  /* fpu.vhdl:1146:57  */
  assign n14711_o = ~n14710_o;
  /* fpu.vhdl:1146:36  */
  assign n14712_o = n14709_o & n14711_o;
  assign n14714_o = r[151];
  /* fpu.vhdl:1146:17  */
  assign n14715_o = n14712_o ? 1'b1 : n14714_o;
  /* fpu.vhdl:1146:17  */
  assign n14718_o = n14712_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1153:24  */
  assign n14720_o = r[318:239];
  /* fpu.vhdl:1153:26  */
  assign n14721_o = n14720_o[1:0];
  /* fpu.vhdl:1154:21  */
  assign n14723_o = n14721_o == 2'b00;
  /* fpu.vhdl:1157:30  */
  assign n14724_o = r[318:239];
  /* fpu.vhdl:1157:32  */
  assign n14725_o = n14724_o[15:3];
  /* fpu.vhdl:1157:41  */
  assign n14727_o = $signed(n14725_o) >= $signed(13'b0000001000000);
  /* fpu.vhdl:1158:36  */
  assign n14728_o = r[26];
  /* fpu.vhdl:1158:40  */
  assign n14729_o = ~n14728_o;
  /* fpu.vhdl:1158:52  */
  assign n14730_o = r[318:239];
  /* fpu.vhdl:1158:54  */
  assign n14731_o = n14730_o[15:3];
  /* fpu.vhdl:1158:63  */
  assign n14733_o = $signed(n14731_o) >= $signed(13'b0000000100000);
  /* fpu.vhdl:1158:46  */
  assign n14734_o = n14729_o & n14733_o;
  /* fpu.vhdl:1157:68  */
  assign n14735_o = n14727_o | n14734_o;
  /* fpu.vhdl:1160:33  */
  assign n14737_o = r[318:239];
  /* fpu.vhdl:1160:35  */
  assign n14738_o = n14737_o[15:3];
  /* fpu.vhdl:1160:44  */
  assign n14740_o = $signed(n14738_o) >= $signed(13'b0000000110100);
  /* fpu.vhdl:1163:42  */
  assign n14741_o = r[318:239];
  /* fpu.vhdl:1163:44  */
  assign n14742_o = n14741_o[15:3];
  /* fpu.vhdl:1163:53  */
  assign n14744_o = n14742_o - 13'b0000000110110;
  /* fpu.vhdl:1164:38  */
  assign n14745_o = r[25];
  /* fpu.vhdl:1164:54  */
  assign n14746_o = r[318:239];
  /* fpu.vhdl:1164:56  */
  assign n14747_o = n14746_o[2];
  /* fpu.vhdl:1164:48  */
  assign n14748_o = n14745_o & n14747_o;
  /* fpu.vhdl:1164:29  */
  assign n14751_o = n14748_o ? 7'b0111111 : 7'b0111100;
  /* fpu.vhdl:1170:42  */
  assign n14752_o = r[318:239];
  /* fpu.vhdl:1170:44  */
  assign n14753_o = n14752_o[15:3];
  /* fpu.vhdl:1170:53  */
  assign n14755_o = n14753_o - 13'b0000000110100;
  /* fpu.vhdl:1160:25  */
  assign n14757_o = n14740_o ? n14751_o : 7'b0111010;
  /* fpu.vhdl:1160:25  */
  assign n14758_o = n14740_o ? n14744_o : n14755_o;
  /* fpu.vhdl:1157:25  */
  assign n14759_o = n14735_o ? 7'b0111111 : n14757_o;
  /* fpu.vhdl:1157:25  */
  assign n14760_o = n14735_o ? 13'b0000000000000 : n14758_o;
  /* fpu.vhdl:1156:21  */
  assign n14762_o = n14721_o == 2'b01;
  /* fpu.vhdl:1173:21  */
  assign n14765_o = n14721_o == 2'b10;
  /* fpu.vhdl:1173:35  */
  assign n14767_o = n14721_o == 2'b11;
  /* fpu.vhdl:1173:35  */
  assign n14768_o = n14765_o | n14767_o;
  assign n14769_o = {n14768_o, n14762_o, n14723_o};
  /* fpu.vhdl:1153:17  */
  always @*
    case (n14769_o)
      3'b100: n14771_o = 7'b0111111;
      3'b010: n14771_o = n14759_o;
      3'b001: n14771_o = n13151_o;
      default: n14771_o = 7'bX;
    endcase
  /* fpu.vhdl:1153:17  */
  always @*
    case (n14769_o)
      3'b100: n14773_o = 13'b0000000000000;
      3'b010: n14773_o = n14760_o;
      3'b001: n14773_o = 13'b0000000000000;
      default: n14773_o = 13'bX;
    endcase
  /* fpu.vhdl:1153:17  */
  always @*
    case (n14769_o)
      3'b100: n14777_o = 1'b0;
      3'b010: n14777_o = 1'b0;
      3'b001: n14777_o = 1'b1;
      default: n14777_o = 1'bX;
    endcase
  /* fpu.vhdl:1136:13  */
  assign n14779_o = n13567_o == 7'b0001100;
  /* fpu.vhdl:1180:26  */
  assign n14781_o = r[25];
  /* fpu.vhdl:1180:30  */
  assign n14782_o = ~n14781_o;
  /* fpu.vhdl:1180:42  */
  assign n14783_o = r[318:239];
  /* fpu.vhdl:1180:44  */
  assign n14784_o = n14783_o[2];
  /* fpu.vhdl:1180:36  */
  assign n14785_o = n14782_o & n14784_o;
  /* fpu.vhdl:1180:17  */
  assign n14789_o = n14785_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1180:17  */
  assign n14792_o = n14785_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1180:17  */
  assign n14793_o = n14785_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1186:37  */
  assign n14794_o = r[318:239];
  /* fpu.vhdl:1186:39  */
  assign n14795_o = n14794_o[1:0];
  /* fpu.vhdl:1190:22  */
  assign n14799_o = r[318:239];
  /* fpu.vhdl:1190:24  */
  assign n14800_o = n14799_o[1:0];
  /* fpu.vhdl:1190:30  */
  assign n14802_o = n14800_o == 2'b00;
  /* fpu.vhdl:1190:17  */
  assign n14804_o = n14802_o ? n13151_o : 7'b1000000;
  /* fpu.vhdl:1190:17  */
  assign n14807_o = n14802_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1177:13  */
  assign n14809_o = n13567_o == 7'b0001011;
  /* fpu.vhdl:1199:36  */
  assign n14810_o = r[238:159];
  /* fpu.vhdl:1199:38  */
  assign n14811_o = n14810_o[2];
  /* fpu.vhdl:1200:37  */
  assign n14812_o = r[238:159];
  /* fpu.vhdl:1200:39  */
  assign n14813_o = n14812_o[1:0];
  /* fpu.vhdl:1201:35  */
  assign n14814_o = r[238:159];
  /* fpu.vhdl:1201:37  */
  assign n14815_o = n14814_o[15:3];
  /* fpu.vhdl:1206:29  */
  assign n14820_o = r[238:159];
  /* fpu.vhdl:1206:31  */
  assign n14821_o = n14820_o[2];
  /* fpu.vhdl:1206:46  */
  assign n14822_o = r[318:239];
  /* fpu.vhdl:1206:48  */
  assign n14823_o = n14822_o[2];
  /* fpu.vhdl:1206:40  */
  assign n14824_o = n14821_o ^ n14823_o;
  /* fpu.vhdl:1206:67  */
  assign n14825_o = r[18];
  /* fpu.vhdl:1206:57  */
  assign n14826_o = n14824_o ^ n14825_o;
  /* fpu.vhdl:1207:22  */
  assign n14827_o = r[238:159];
  /* fpu.vhdl:1207:24  */
  assign n14828_o = n14827_o[1:0];
  /* fpu.vhdl:1207:30  */
  assign n14830_o = n14828_o == 2'b01;
  /* fpu.vhdl:1207:45  */
  assign n14831_o = r[318:239];
  /* fpu.vhdl:1207:47  */
  assign n14832_o = n14831_o[1:0];
  /* fpu.vhdl:1207:53  */
  assign n14834_o = n14832_o == 2'b01;
  /* fpu.vhdl:1207:39  */
  assign n14835_o = n14830_o & n14834_o;
  /* fpu.vhdl:1208:38  */
  assign n14836_o = ~n14826_o;
  /* fpu.vhdl:1209:39  */
  assign n14837_o = r[704];
  /* fpu.vhdl:1211:26  */
  assign n14839_o = r[704];
  /* fpu.vhdl:1211:34  */
  assign n14840_o = ~n14839_o;
  /* fpu.vhdl:1212:38  */
  assign n14841_o = r[238:159];
  /* fpu.vhdl:1212:40  */
  assign n14842_o = n14841_o[15:3];
  /* fpu.vhdl:1212:53  */
  assign n14843_o = r[318:239];
  /* fpu.vhdl:1212:55  */
  assign n14844_o = n14843_o[15:3];
  /* fpu.vhdl:1212:49  */
  assign n14845_o = n14842_o - n14844_o;
  /* fpu.vhdl:1213:44  */
  assign n14846_o = r[318:239];
  /* fpu.vhdl:1213:46  */
  assign n14847_o = n14846_o[2];
  /* fpu.vhdl:1213:66  */
  assign n14848_o = r[18];
  /* fpu.vhdl:1213:55  */
  assign n14849_o = ~(n14847_o ^ n14848_o);
  /* fpu.vhdl:1214:30  */
  assign n14850_o = r[238:159];
  /* fpu.vhdl:1214:32  */
  assign n14851_o = n14850_o[15:3];
  /* fpu.vhdl:1214:45  */
  assign n14852_o = r[318:239];
  /* fpu.vhdl:1214:47  */
  assign n14853_o = n14852_o[15:3];
  /* fpu.vhdl:1214:41  */
  assign n14854_o = n14851_o == n14853_o;
  /* fpu.vhdl:1214:25  */
  assign n14858_o = n14854_o ? 7'b0011010 : 7'b0011001;
  /* fpu.vhdl:1214:25  */
  assign n14859_o = n14854_o ? n13479_o : 1'b0;
  /* fpu.vhdl:1211:21  */
  assign n14861_o = n14840_o ? n14858_o : 7'b0011000;
  /* fpu.vhdl:1211:21  */
  assign n14862_o = n14840_o ? n14849_o : n14811_o;
  /* fpu.vhdl:1207:17  */
  assign n14863_o = n14955_o ? n14845_o : 13'b0000000000000;
  /* fpu.vhdl:1207:17  */
  assign n14864_o = n14967_o ? n14859_o : n13479_o;
  /* fpu.vhdl:1224:26  */
  assign n14865_o = r[238:159];
  /* fpu.vhdl:1224:28  */
  assign n14866_o = n14865_o[1:0];
  /* fpu.vhdl:1224:34  */
  assign n14868_o = n14866_o == 2'b11;
  /* fpu.vhdl:1224:45  */
  assign n14869_o = r[318:239];
  /* fpu.vhdl:1224:47  */
  assign n14870_o = n14869_o[1:0];
  /* fpu.vhdl:1224:53  */
  assign n14872_o = n14870_o == 2'b11;
  /* fpu.vhdl:1224:40  */
  assign n14873_o = n14868_o | n14872_o;
  /* fpu.vhdl:1226:29  */
  assign n14875_o = r[238:159];
  /* fpu.vhdl:1226:31  */
  assign n14876_o = n14875_o[1:0];
  /* fpu.vhdl:1226:37  */
  assign n14878_o = n14876_o == 2'b10;
  /* fpu.vhdl:1226:54  */
  assign n14879_o = r[318:239];
  /* fpu.vhdl:1226:56  */
  assign n14880_o = n14879_o[1:0];
  /* fpu.vhdl:1226:62  */
  assign n14882_o = n14880_o == 2'b10;
  /* fpu.vhdl:1226:48  */
  assign n14883_o = n14878_o & n14882_o;
  /* fpu.vhdl:1226:84  */
  assign n14884_o = ~n14826_o;
  /* fpu.vhdl:1226:73  */
  assign n14885_o = n14883_o & n14884_o;
  /* fpu.vhdl:1231:29  */
  assign n14887_o = r[238:159];
  /* fpu.vhdl:1231:31  */
  assign n14888_o = n14887_o[1:0];
  /* fpu.vhdl:1231:37  */
  assign n14890_o = n14888_o == 2'b00;
  /* fpu.vhdl:1231:50  */
  assign n14891_o = r[318:239];
  /* fpu.vhdl:1231:52  */
  assign n14892_o = n14891_o[1:0];
  /* fpu.vhdl:1231:58  */
  assign n14894_o = n14892_o == 2'b00;
  /* fpu.vhdl:1231:44  */
  assign n14895_o = n14890_o & n14894_o;
  /* fpu.vhdl:1231:76  */
  assign n14896_o = ~n14826_o;
  /* fpu.vhdl:1231:65  */
  assign n14897_o = n14895_o & n14896_o;
  /* fpu.vhdl:1233:54  */
  assign n14898_o = r[701];
  /* fpu.vhdl:1233:74  */
  assign n14899_o = r[700];
  /* fpu.vhdl:1233:58  */
  assign n14900_o = n14898_o & n14899_o;
  /* fpu.vhdl:1235:29  */
  assign n14901_o = r[238:159];
  /* fpu.vhdl:1235:31  */
  assign n14902_o = n14901_o[1:0];
  /* fpu.vhdl:1235:37  */
  assign n14904_o = n14902_o == 2'b10;
  /* fpu.vhdl:1235:53  */
  assign n14905_o = r[318:239];
  /* fpu.vhdl:1235:55  */
  assign n14906_o = n14905_o[1:0];
  /* fpu.vhdl:1235:61  */
  assign n14908_o = n14906_o == 2'b00;
  /* fpu.vhdl:1235:48  */
  assign n14909_o = n14904_o | n14908_o;
  /* fpu.vhdl:1242:47  */
  assign n14913_o = r[18];
  /* fpu.vhdl:1242:37  */
  assign n14914_o = ~n14913_o;
  /* fpu.vhdl:1235:21  */
  assign n14916_o = n14909_o ? 7'b1001111 : 7'b1001111;
  /* fpu.vhdl:1235:21  */
  assign n14917_o = n14909_o ? 2'b01 : 2'b10;
  assign n14918_o = r[720];
  /* fpu.vhdl:1235:21  */
  assign n14919_o = n14909_o ? n14918_o : n14914_o;
  /* fpu.vhdl:1231:21  */
  assign n14920_o = n14897_o ? n13151_o : n14916_o;
  /* fpu.vhdl:1231:21  */
  assign n14921_o = n14897_o ? n14900_o : n14811_o;
  /* fpu.vhdl:1231:21  */
  assign n14922_o = n14897_o ? 2'b00 : n14917_o;
  assign n14923_o = r[720];
  /* fpu.vhdl:1231:21  */
  assign n14924_o = n14897_o ? n14923_o : n14919_o;
  /* fpu.vhdl:1231:21  */
  assign n14927_o = n14897_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1226:21  */
  assign n14928_o = n14885_o ? n13151_o : n14920_o;
  assign n14929_o = r[150];
  /* fpu.vhdl:1226:21  */
  assign n14930_o = n14885_o ? 1'b1 : n14929_o;
  /* fpu.vhdl:1226:21  */
  assign n14931_o = n14885_o ? n14811_o : n14921_o;
  /* fpu.vhdl:1226:21  */
  assign n14932_o = n14885_o ? 2'b00 : n14922_o;
  assign n14933_o = r[720];
  /* fpu.vhdl:1226:21  */
  assign n14934_o = n14885_o ? n14933_o : n14924_o;
  /* fpu.vhdl:1226:21  */
  assign n14936_o = n14885_o ? 1'b1 : n14927_o;
  /* fpu.vhdl:1226:21  */
  assign n14939_o = n14885_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1224:21  */
  assign n14940_o = n14873_o ? 7'b1001110 : n14928_o;
  assign n14941_o = r[150];
  /* fpu.vhdl:1224:21  */
  assign n14942_o = n14873_o ? n14941_o : n14930_o;
  /* fpu.vhdl:1224:21  */
  assign n14943_o = n14873_o ? n14811_o : n14931_o;
  /* fpu.vhdl:1224:21  */
  assign n14944_o = n14873_o ? 2'b00 : n14932_o;
  assign n14945_o = r[720];
  /* fpu.vhdl:1224:21  */
  assign n14946_o = n14873_o ? n14945_o : n14934_o;
  /* fpu.vhdl:1224:21  */
  assign n14948_o = n14873_o ? 1'b0 : n14936_o;
  /* fpu.vhdl:1224:21  */
  assign n14950_o = n14873_o ? 1'b0 : n14939_o;
  /* fpu.vhdl:1207:17  */
  assign n14951_o = n14835_o ? n14861_o : n14940_o;
  assign n14952_o = r[150];
  /* fpu.vhdl:1207:17  */
  assign n14953_o = n14835_o ? n14952_o : n14942_o;
  /* fpu.vhdl:1207:17  */
  assign n14954_o = n14835_o ? n14862_o : n14943_o;
  /* fpu.vhdl:1207:17  */
  assign n14955_o = n14835_o & n14840_o;
  assign n14956_o = n13465_o[6];
  assign n14957_o = r[703];
  /* fpu.vhdl:650:9  */
  assign n14958_o = n13152_o ? n14956_o : n14957_o;
  /* fpu.vhdl:1207:17  */
  assign n14959_o = n14835_o ? n14836_o : n14958_o;
  assign n14960_o = n13465_o[9];
  assign n14961_o = r[706];
  /* fpu.vhdl:650:9  */
  assign n14962_o = n13152_o ? n14960_o : n14961_o;
  /* fpu.vhdl:1207:17  */
  assign n14963_o = n14835_o ? n14837_o : n14962_o;
  /* fpu.vhdl:1207:17  */
  assign n14964_o = n14835_o ? 2'b10 : n14944_o;
  assign n14965_o = r[720];
  /* fpu.vhdl:1207:17  */
  assign n14966_o = n14835_o ? n14965_o : n14946_o;
  /* fpu.vhdl:1207:17  */
  assign n14967_o = n14835_o & n14840_o;
  /* fpu.vhdl:1207:17  */
  assign n14969_o = n14835_o ? 1'b0 : n14948_o;
  /* fpu.vhdl:1207:17  */
  assign n14971_o = n14835_o ? 1'b0 : n14950_o;
  /* fpu.vhdl:1196:13  */
  assign n14973_o = n13567_o == 7'b0001111;
  /* fpu.vhdl:1250:36  */
  assign n14974_o = r[238:159];
  /* fpu.vhdl:1250:38  */
  assign n14975_o = n14974_o[2];
  /* fpu.vhdl:1250:53  */
  assign n14976_o = r[398:319];
  /* fpu.vhdl:1250:55  */
  assign n14977_o = n14976_o[2];
  /* fpu.vhdl:1250:47  */
  assign n14978_o = n14975_o ^ n14977_o;
  /* fpu.vhdl:1251:37  */
  assign n14979_o = r[238:159];
  /* fpu.vhdl:1251:39  */
  assign n14980_o = n14979_o[1:0];
  /* fpu.vhdl:1256:22  */
  assign n14985_o = r[238:159];
  /* fpu.vhdl:1256:24  */
  assign n14986_o = n14985_o[1:0];
  /* fpu.vhdl:1256:30  */
  assign n14988_o = n14986_o == 2'b01;
  /* fpu.vhdl:1256:45  */
  assign n14989_o = r[398:319];
  /* fpu.vhdl:1256:47  */
  assign n14990_o = n14989_o[1:0];
  /* fpu.vhdl:1256:53  */
  assign n14992_o = n14990_o == 2'b01;
  /* fpu.vhdl:1256:39  */
  assign n14993_o = n14988_o & n14992_o;
  /* fpu.vhdl:1257:39  */
  assign n14994_o = r[238:159];
  /* fpu.vhdl:1257:41  */
  assign n14995_o = n14994_o[15:3];
  /* fpu.vhdl:1257:54  */
  assign n14996_o = r[398:319];
  /* fpu.vhdl:1257:56  */
  assign n14997_o = n14996_o[15:3];
  /* fpu.vhdl:1257:50  */
  assign n14998_o = n14995_o + n14997_o;
  /* fpu.vhdl:1259:36  */
  assign n14999_o = r[229];
  /* fpu.vhdl:1259:41  */
  assign n15000_o = ~n14999_o;
  /* fpu.vhdl:1261:39  */
  assign n15002_o = r[389];
  /* fpu.vhdl:1261:44  */
  assign n15003_o = ~n15002_o;
  /* fpu.vhdl:1261:21  */
  assign n15007_o = n15003_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:1261:21  */
  assign n15008_o = n15003_o ? 7'b1001100 : 7'b0011110;
  /* fpu.vhdl:1259:21  */
  assign n15009_o = n15000_o ? 1'b0 : n15007_o;
  /* fpu.vhdl:1259:21  */
  assign n15010_o = n15000_o ? 7'b1001000 : n15008_o;
  /* fpu.vhdl:1268:26  */
  assign n15011_o = r[238:159];
  /* fpu.vhdl:1268:28  */
  assign n15012_o = n15011_o[1:0];
  /* fpu.vhdl:1268:34  */
  assign n15014_o = n15012_o == 2'b11;
  /* fpu.vhdl:1268:45  */
  assign n15015_o = r[398:319];
  /* fpu.vhdl:1268:47  */
  assign n15016_o = n15015_o[1:0];
  /* fpu.vhdl:1268:53  */
  assign n15018_o = n15016_o == 2'b11;
  /* fpu.vhdl:1268:40  */
  assign n15019_o = n15014_o | n15018_o;
  /* fpu.vhdl:1270:30  */
  assign n15021_o = r[238:159];
  /* fpu.vhdl:1270:32  */
  assign n15022_o = n15021_o[1:0];
  /* fpu.vhdl:1270:38  */
  assign n15024_o = n15022_o == 2'b10;
  /* fpu.vhdl:1270:55  */
  assign n15025_o = r[398:319];
  /* fpu.vhdl:1270:57  */
  assign n15026_o = n15025_o[1:0];
  /* fpu.vhdl:1270:63  */
  assign n15028_o = n15026_o == 2'b00;
  /* fpu.vhdl:1270:49  */
  assign n15029_o = n15024_o & n15028_o;
  /* fpu.vhdl:1271:28  */
  assign n15030_o = r[238:159];
  /* fpu.vhdl:1271:30  */
  assign n15031_o = n15030_o[1:0];
  /* fpu.vhdl:1271:36  */
  assign n15033_o = n15031_o == 2'b00;
  /* fpu.vhdl:1271:49  */
  assign n15034_o = r[398:319];
  /* fpu.vhdl:1271:51  */
  assign n15035_o = n15034_o[1:0];
  /* fpu.vhdl:1271:57  */
  assign n15037_o = n15035_o == 2'b10;
  /* fpu.vhdl:1271:43  */
  assign n15038_o = n15033_o & n15037_o;
  /* fpu.vhdl:1270:71  */
  assign n15039_o = n15029_o | n15038_o;
  /* fpu.vhdl:1275:29  */
  assign n15041_o = r[238:159];
  /* fpu.vhdl:1275:31  */
  assign n15042_o = n15041_o[1:0];
  /* fpu.vhdl:1275:37  */
  assign n15044_o = n15042_o == 2'b00;
  /* fpu.vhdl:1275:49  */
  assign n15045_o = r[238:159];
  /* fpu.vhdl:1275:51  */
  assign n15046_o = n15045_o[1:0];
  /* fpu.vhdl:1275:57  */
  assign n15048_o = n15046_o == 2'b10;
  /* fpu.vhdl:1275:44  */
  assign n15049_o = n15044_o | n15048_o;
  /* fpu.vhdl:1281:39  */
  assign n15051_o = r[238:159];
  /* fpu.vhdl:1281:41  */
  assign n15052_o = n15051_o[2];
  /* fpu.vhdl:1275:21  */
  assign n15054_o = n15049_o ? n13151_o : 7'b1001111;
  /* fpu.vhdl:1275:21  */
  assign n15055_o = n15049_o ? 2'b00 : 2'b11;
  assign n15056_o = r[720];
  /* fpu.vhdl:1275:21  */
  assign n15057_o = n15049_o ? n15056_o : n15052_o;
  /* fpu.vhdl:1275:21  */
  assign n15060_o = n15049_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1270:21  */
  assign n15061_o = n15039_o ? n13151_o : n15054_o;
  assign n15062_o = r[147];
  /* fpu.vhdl:1270:21  */
  assign n15063_o = n15039_o ? 1'b1 : n15062_o;
  /* fpu.vhdl:1270:21  */
  assign n15064_o = n15039_o ? 2'b00 : n15055_o;
  assign n15065_o = r[720];
  /* fpu.vhdl:1270:21  */
  assign n15066_o = n15039_o ? n15065_o : n15057_o;
  /* fpu.vhdl:1270:21  */
  assign n15068_o = n15039_o ? 1'b0 : n15060_o;
  /* fpu.vhdl:1270:21  */
  assign n15071_o = n15039_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1268:21  */
  assign n15072_o = n15019_o ? 7'b1001110 : n15061_o;
  assign n15073_o = r[147];
  /* fpu.vhdl:1268:21  */
  assign n15074_o = n15019_o ? n15073_o : n15063_o;
  /* fpu.vhdl:1268:21  */
  assign n15075_o = n15019_o ? 2'b00 : n15064_o;
  assign n15076_o = r[720];
  /* fpu.vhdl:1268:21  */
  assign n15077_o = n15019_o ? n15076_o : n15066_o;
  /* fpu.vhdl:1268:21  */
  assign n15079_o = n15019_o ? 1'b0 : n15068_o;
  /* fpu.vhdl:1268:21  */
  assign n15081_o = n15019_o ? 1'b0 : n15071_o;
  /* fpu.vhdl:1256:17  */
  assign n15082_o = n14993_o ? n15009_o : 1'b0;
  /* fpu.vhdl:1256:17  */
  assign n15083_o = n14993_o ? n15010_o : n15072_o;
  assign n15084_o = r[147];
  /* fpu.vhdl:1256:17  */
  assign n15085_o = n14993_o ? n15084_o : n15074_o;
  assign n15086_o = r[663:651];
  /* fpu.vhdl:1256:17  */
  assign n15087_o = n14993_o ? n14998_o : n15086_o;
  /* fpu.vhdl:1256:17  */
  assign n15088_o = n14993_o ? 2'b00 : n15075_o;
  assign n15089_o = r[720];
  /* fpu.vhdl:1256:17  */
  assign n15090_o = n14993_o ? n15089_o : n15077_o;
  /* fpu.vhdl:1256:17  */
  assign n15092_o = n14993_o ? 1'b0 : n15079_o;
  /* fpu.vhdl:1256:17  */
  assign n15094_o = n14993_o ? 1'b0 : n15081_o;
  /* fpu.vhdl:1247:13  */
  assign n15096_o = n13567_o == 7'b0010000;
  /* fpu.vhdl:1288:37  */
  assign n15097_o = r[238:159];
  /* fpu.vhdl:1288:39  */
  assign n15098_o = n15097_o[1:0];
  /* fpu.vhdl:1293:36  */
  assign n15103_o = r[238:159];
  /* fpu.vhdl:1293:38  */
  assign n15104_o = n15103_o[2];
  /* fpu.vhdl:1293:53  */
  assign n15105_o = r[318:239];
  /* fpu.vhdl:1293:55  */
  assign n15106_o = n15105_o[2];
  /* fpu.vhdl:1293:47  */
  assign n15107_o = n15104_o ^ n15106_o;
  /* fpu.vhdl:1294:35  */
  assign n15108_o = r[238:159];
  /* fpu.vhdl:1294:37  */
  assign n15109_o = n15108_o[15:3];
  /* fpu.vhdl:1294:50  */
  assign n15110_o = r[318:239];
  /* fpu.vhdl:1294:52  */
  assign n15111_o = n15110_o[15:3];
  /* fpu.vhdl:1294:46  */
  assign n15112_o = n15109_o - n15111_o;
  /* fpu.vhdl:1296:22  */
  assign n15114_o = r[238:159];
  /* fpu.vhdl:1296:24  */
  assign n15115_o = n15114_o[1:0];
  /* fpu.vhdl:1296:30  */
  assign n15117_o = n15115_o == 2'b01;
  /* fpu.vhdl:1296:45  */
  assign n15118_o = r[318:239];
  /* fpu.vhdl:1296:47  */
  assign n15119_o = n15118_o[1:0];
  /* fpu.vhdl:1296:53  */
  assign n15121_o = n15119_o == 2'b01;
  /* fpu.vhdl:1296:39  */
  assign n15122_o = n15117_o & n15121_o;
  /* fpu.vhdl:1298:36  */
  assign n15123_o = r[229];
  /* fpu.vhdl:1298:41  */
  assign n15124_o = ~n15123_o;
  /* fpu.vhdl:1300:39  */
  assign n15126_o = r[309];
  /* fpu.vhdl:1300:44  */
  assign n15127_o = ~n15126_o;
  /* fpu.vhdl:1300:21  */
  assign n15131_o = n15127_o ? 7'b1001010 : 7'b0100110;
  /* fpu.vhdl:1300:21  */
  assign n15132_o = n15127_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:1298:21  */
  assign n15133_o = n15124_o ? 7'b1001000 : n15131_o;
  /* fpu.vhdl:1298:21  */
  assign n15134_o = n15124_o ? 1'b0 : n15132_o;
  /* fpu.vhdl:1307:26  */
  assign n15135_o = r[238:159];
  /* fpu.vhdl:1307:28  */
  assign n15136_o = n15135_o[1:0];
  /* fpu.vhdl:1307:34  */
  assign n15138_o = n15136_o == 2'b11;
  /* fpu.vhdl:1307:45  */
  assign n15139_o = r[318:239];
  /* fpu.vhdl:1307:47  */
  assign n15140_o = n15139_o[1:0];
  /* fpu.vhdl:1307:53  */
  assign n15142_o = n15140_o == 2'b11;
  /* fpu.vhdl:1307:40  */
  assign n15143_o = n15138_o | n15142_o;
  /* fpu.vhdl:1309:29  */
  assign n15145_o = r[318:239];
  /* fpu.vhdl:1309:31  */
  assign n15146_o = n15145_o[1:0];
  /* fpu.vhdl:1309:37  */
  assign n15148_o = n15146_o == 2'b10;
  /* fpu.vhdl:1310:30  */
  assign n15149_o = r[238:159];
  /* fpu.vhdl:1310:32  */
  assign n15150_o = n15149_o[1:0];
  /* fpu.vhdl:1310:38  */
  assign n15152_o = n15150_o == 2'b10;
  assign n15155_o = r[149];
  /* fpu.vhdl:1309:21  */
  assign n15156_o = n15196_o ? 1'b1 : n15155_o;
  /* fpu.vhdl:1310:25  */
  assign n15157_o = n15152_o ? n15098_o : 2'b00;
  /* fpu.vhdl:1310:25  */
  assign n15160_o = n15152_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1317:29  */
  assign n15161_o = r[318:239];
  /* fpu.vhdl:1317:31  */
  assign n15162_o = n15161_o[1:0];
  /* fpu.vhdl:1317:37  */
  assign n15164_o = n15162_o == 2'b00;
  /* fpu.vhdl:1318:30  */
  assign n15165_o = r[238:159];
  /* fpu.vhdl:1318:32  */
  assign n15166_o = n15165_o[1:0];
  /* fpu.vhdl:1318:38  */
  assign n15168_o = n15166_o == 2'b00;
  /* fpu.vhdl:1322:34  */
  assign n15170_o = r[238:159];
  /* fpu.vhdl:1322:36  */
  assign n15171_o = n15170_o[1:0];
  /* fpu.vhdl:1322:42  */
  assign n15173_o = n15171_o == 2'b01;
  /* fpu.vhdl:1322:29  */
  assign n15176_o = n15173_o ? 1'b1 : 1'b0;
  assign n15178_o = r[148];
  /* fpu.vhdl:1317:21  */
  assign n15179_o = n15187_o ? 1'b1 : n15178_o;
  /* fpu.vhdl:1318:25  */
  assign n15180_o = n15168_o ? n15098_o : 2'b10;
  /* fpu.vhdl:1318:25  */
  assign n15182_o = n15168_o ? 1'b0 : n15176_o;
  /* fpu.vhdl:1318:25  */
  assign n15185_o = n15168_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1317:21  */
  assign n15187_o = n15164_o & n15168_o;
  /* fpu.vhdl:1317:21  */
  assign n15188_o = n15164_o ? n15180_o : n15098_o;
  /* fpu.vhdl:1317:21  */
  assign n15190_o = n15164_o ? n15182_o : 1'b0;
  /* fpu.vhdl:1317:21  */
  assign n15192_o = n15164_o ? n15185_o : 1'b0;
  assign n15193_o = r[148];
  /* fpu.vhdl:1309:21  */
  assign n15194_o = n15148_o ? n15193_o : n15179_o;
  /* fpu.vhdl:1309:21  */
  assign n15196_o = n15148_o & n15152_o;
  /* fpu.vhdl:1309:21  */
  assign n15197_o = n15148_o ? n15157_o : n15188_o;
  /* fpu.vhdl:1309:21  */
  assign n15199_o = n15148_o ? 1'b0 : n15190_o;
  /* fpu.vhdl:1309:21  */
  assign n15200_o = n15148_o ? n15160_o : n15192_o;
  assign n15201_o = {n15156_o, n15194_o};
  /* fpu.vhdl:1307:21  */
  assign n15202_o = n15143_o ? 7'b1001110 : n13151_o;
  assign n15203_o = r[149:148];
  /* fpu.vhdl:1307:21  */
  assign n15204_o = n15143_o ? n15203_o : n15201_o;
  /* fpu.vhdl:1307:21  */
  assign n15205_o = n15143_o ? n15098_o : n15197_o;
  /* fpu.vhdl:1307:21  */
  assign n15208_o = n15143_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:1307:21  */
  assign n15210_o = n15143_o ? 1'b0 : n15199_o;
  /* fpu.vhdl:1307:21  */
  assign n15212_o = n15143_o ? 1'b0 : n15200_o;
  /* fpu.vhdl:1296:17  */
  assign n15213_o = n15122_o ? n15133_o : n15202_o;
  assign n15214_o = r[149:148];
  /* fpu.vhdl:1296:17  */
  assign n15215_o = n15122_o ? n15214_o : n15204_o;
  /* fpu.vhdl:1296:17  */
  assign n15216_o = n15122_o ? n15098_o : n15205_o;
  /* fpu.vhdl:1296:17  */
  assign n15217_o = n15122_o ? n15134_o : 1'b0;
  /* fpu.vhdl:1296:17  */
  assign n15219_o = n15122_o ? 1'b0 : n15208_o;
  /* fpu.vhdl:1296:17  */
  assign n15221_o = n15122_o ? 1'b0 : n15210_o;
  /* fpu.vhdl:1296:17  */
  assign n15223_o = n15122_o ? 1'b0 : n15212_o;
  /* fpu.vhdl:1286:13  */
  assign n15225_o = n13567_o == 7'b0010001;
  /* fpu.vhdl:1336:22  */
  assign n15228_o = r[238:159];
  /* fpu.vhdl:1336:24  */
  assign n15229_o = n15228_o[1:0];
  /* fpu.vhdl:1336:30  */
  assign n15231_o = n15229_o == 2'b00;
  /* fpu.vhdl:1336:43  */
  assign n15232_o = r[238:159];
  /* fpu.vhdl:1336:45  */
  assign n15233_o = n15232_o[2];
  /* fpu.vhdl:1336:54  */
  assign n15234_o = ~n15233_o;
  /* fpu.vhdl:1336:66  */
  assign n15235_o = r[238:159];
  /* fpu.vhdl:1336:68  */
  assign n15236_o = n15235_o[1:0];
  /* fpu.vhdl:1336:74  */
  assign n15238_o = n15236_o != 2'b11;
  /* fpu.vhdl:1336:60  */
  assign n15239_o = n15234_o & n15238_o;
  /* fpu.vhdl:1336:37  */
  assign n15240_o = n15231_o | n15239_o;
  /* fpu.vhdl:1336:17  */
  assign n15243_o = n15240_o ? 2'b11 : 2'b10;
  /* fpu.vhdl:1333:13  */
  assign n15247_o = n13567_o == 7'b0010110;
  /* fpu.vhdl:1346:37  */
  assign n15248_o = r[318:239];
  /* fpu.vhdl:1346:39  */
  assign n15249_o = n15248_o[1:0];
  /* fpu.vhdl:1347:36  */
  assign n15250_o = r[318:239];
  /* fpu.vhdl:1347:38  */
  assign n15251_o = n15250_o[2];
  /* fpu.vhdl:1351:24  */
  assign n15255_o = r[318:239];
  /* fpu.vhdl:1351:26  */
  assign n15256_o = n15255_o[1:0];
  /* fpu.vhdl:1353:43  */
  assign n15257_o = r[318:239];
  /* fpu.vhdl:1353:45  */
  assign n15258_o = n15257_o[15:3];
  /* fpu.vhdl:1354:30  */
  assign n15259_o = r[318:239];
  /* fpu.vhdl:1354:32  */
  assign n15260_o = n15259_o[2];
  /* fpu.vhdl:1357:43  */
  assign n15262_o = r[309];
  /* fpu.vhdl:1357:48  */
  assign n15263_o = ~n15262_o;
  /* fpu.vhdl:1359:43  */
  assign n15265_o = r[242];
  /* fpu.vhdl:1359:47  */
  assign n15266_o = ~n15265_o;
  /* fpu.vhdl:1359:25  */
  assign n15270_o = n15266_o ? 7'b0101110 : 7'b1001011;
  /* fpu.vhdl:1359:25  */
  assign n15271_o = n15266_o ? 13'b0000000000000 : 13'b0000000000001;
  /* fpu.vhdl:1357:25  */
  assign n15272_o = n15263_o ? 7'b1001010 : n15270_o;
  /* fpu.vhdl:1357:25  */
  assign n15273_o = n15263_o ? 13'b0000000000000 : n15271_o;
  /* fpu.vhdl:1354:25  */
  assign n15274_o = n15260_o ? n13151_o : n15272_o;
  assign n15275_o = r[136];
  /* fpu.vhdl:1354:25  */
  assign n15276_o = n15260_o ? 1'b1 : n15275_o;
  /* fpu.vhdl:1354:25  */
  assign n15277_o = n15260_o ? 13'b0000000000000 : n15273_o;
  /* fpu.vhdl:1354:25  */
  assign n15280_o = n15260_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1352:21  */
  assign n15282_o = n15256_o == 2'b01;
  /* fpu.vhdl:1365:21  */
  assign n15285_o = n15256_o == 2'b11;
  /* fpu.vhdl:1367:21  */
  assign n15287_o = n15256_o == 2'b00;
  /* fpu.vhdl:1371:30  */
  assign n15288_o = r[318:239];
  /* fpu.vhdl:1371:32  */
  assign n15289_o = n15288_o[2];
  assign n15291_o = r[136];
  /* fpu.vhdl:1371:25  */
  assign n15292_o = n15289_o ? 1'b1 : n15291_o;
  /* fpu.vhdl:1371:25  */
  assign n15295_o = n15289_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1370:21  */
  assign n15297_o = n15256_o == 2'b10;
  assign n15298_o = {n15297_o, n15287_o, n15285_o, n15282_o};
  /* fpu.vhdl:1351:17  */
  always @*
    case (n15298_o)
      4'b1000: n15300_o = n13151_o;
      4'b0100: n15300_o = n13151_o;
      4'b0010: n15300_o = 7'b1001110;
      4'b0001: n15300_o = n15274_o;
      default: n15300_o = 7'bX;
    endcase
  assign n15301_o = r[136];
  /* fpu.vhdl:1351:17  */
  always @*
    case (n15298_o)
      4'b1000: n15303_o = n15292_o;
      4'b0100: n15303_o = n15301_o;
      4'b0010: n15303_o = n15301_o;
      4'b0001: n15303_o = n15276_o;
      default: n15303_o = 1'bX;
    endcase
  assign n15304_o = r[663:651];
  /* fpu.vhdl:1351:17  */
  always @*
    case (n15298_o)
      4'b1000: n15306_o = n15304_o;
      4'b0100: n15306_o = n15304_o;
      4'b0010: n15306_o = n15304_o;
      4'b0001: n15306_o = n15258_o;
      default: n15306_o = 13'bX;
    endcase
  /* fpu.vhdl:1351:17  */
  always @*
    case (n15298_o)
      4'b1000: n15308_o = 13'b0000000000000;
      4'b0100: n15308_o = 13'b0000000000000;
      4'b0010: n15308_o = 13'b0000000000000;
      4'b0001: n15308_o = n15277_o;
      default: n15308_o = 13'bX;
    endcase
  /* fpu.vhdl:1351:17  */
  always @*
    case (n15298_o)
      4'b1000: n15313_o = 1'b1;
      4'b0100: n15313_o = 1'b1;
      4'b0010: n15313_o = 1'b0;
      4'b0001: n15313_o = 1'b0;
      default: n15313_o = 1'bX;
    endcase
  /* fpu.vhdl:1351:17  */
  always @*
    case (n15298_o)
      4'b1000: n15316_o = n15295_o;
      4'b0100: n15316_o = 1'b0;
      4'b0010: n15316_o = 1'b0;
      4'b0001: n15316_o = n15280_o;
      default: n15316_o = 1'bX;
    endcase
  /* fpu.vhdl:1344:13  */
  assign n15318_o = n13567_o == 7'b0010010;
  /* fpu.vhdl:1381:37  */
  assign n15319_o = r[318:239];
  /* fpu.vhdl:1381:39  */
  assign n15320_o = n15319_o[1:0];
  /* fpu.vhdl:1382:36  */
  assign n15321_o = r[318:239];
  /* fpu.vhdl:1382:38  */
  assign n15322_o = n15321_o[2];
  /* fpu.vhdl:1386:24  */
  assign n15326_o = r[318:239];
  /* fpu.vhdl:1386:26  */
  assign n15327_o = n15326_o[1:0];
  /* fpu.vhdl:1388:45  */
  assign n15328_o = r[318:239];
  /* fpu.vhdl:1388:47  */
  assign n15329_o = n15328_o[15:3];
  /* fpu.vhdl:1388:41  */
  assign n15330_o = -n15329_o;
  /* fpu.vhdl:1389:40  */
  assign n15331_o = r[309];
  /* fpu.vhdl:1389:45  */
  assign n15332_o = ~n15331_o;
  /* fpu.vhdl:1389:25  */
  assign n15335_o = n15332_o ? 7'b1001010 : 7'b0101011;
  /* fpu.vhdl:1387:21  */
  assign n15337_o = n15327_o == 2'b01;
  /* fpu.vhdl:1394:21  */
  assign n15340_o = n15327_o == 2'b11;
  /* fpu.vhdl:1396:21  */
  assign n15343_o = n15327_o == 2'b10;
  /* fpu.vhdl:1399:21  */
  assign n15346_o = n15327_o == 2'b00;
  assign n15347_o = {n15346_o, n15343_o, n15340_o, n15337_o};
  /* fpu.vhdl:1386:17  */
  always @*
    case (n15347_o)
      4'b1000: n15349_o = n13151_o;
      4'b0100: n15349_o = n13151_o;
      4'b0010: n15349_o = 7'b1001110;
      4'b0001: n15349_o = n15335_o;
      default: n15349_o = 7'bX;
    endcase
  /* fpu.vhdl:1386:17  */
  always @*
    case (n15347_o)
      4'b1000: n15351_o = 2'b10;
      4'b0100: n15351_o = 2'b00;
      4'b0010: n15351_o = n15320_o;
      4'b0001: n15351_o = n15320_o;
      default: n15351_o = 2'bX;
    endcase
  assign n15352_o = r[663:651];
  /* fpu.vhdl:1386:17  */
  always @*
    case (n15347_o)
      4'b1000: n15354_o = n15352_o;
      4'b0100: n15354_o = n15352_o;
      4'b0010: n15354_o = n15352_o;
      4'b0001: n15354_o = n15330_o;
      default: n15354_o = 13'bX;
    endcase
  /* fpu.vhdl:1386:17  */
  always @*
    case (n15347_o)
      4'b1000: n15359_o = 1'b1;
      4'b0100: n15359_o = 1'b1;
      4'b0010: n15359_o = 1'b0;
      4'b0001: n15359_o = 1'b0;
      default: n15359_o = 1'bX;
    endcase
  /* fpu.vhdl:1386:17  */
  always @*
    case (n15347_o)
      4'b1000: n15363_o = 1'b1;
      4'b0100: n15363_o = 1'b0;
      4'b0010: n15363_o = 1'b0;
      4'b0001: n15363_o = 1'b0;
      default: n15363_o = 1'bX;
    endcase
  /* fpu.vhdl:1379:13  */
  assign n15365_o = n13567_o == 7'b0010100;
  /* fpu.vhdl:1407:37  */
  assign n15366_o = r[318:239];
  /* fpu.vhdl:1407:39  */
  assign n15367_o = n15366_o[1:0];
  /* fpu.vhdl:1408:36  */
  assign n15368_o = r[318:239];
  /* fpu.vhdl:1408:38  */
  assign n15369_o = n15368_o[2];
  /* fpu.vhdl:1413:24  */
  assign n15374_o = r[318:239];
  /* fpu.vhdl:1413:26  */
  assign n15375_o = n15374_o[1:0];
  /* fpu.vhdl:1415:43  */
  assign n15376_o = r[318:239];
  /* fpu.vhdl:1415:45  */
  assign n15377_o = n15376_o[15:3];
  /* fpu.vhdl:1416:30  */
  assign n15378_o = r[318:239];
  /* fpu.vhdl:1416:32  */
  assign n15379_o = n15378_o[2];
  /* fpu.vhdl:1419:43  */
  assign n15381_o = r[309];
  /* fpu.vhdl:1419:48  */
  assign n15382_o = ~n15381_o;
  /* fpu.vhdl:1421:43  */
  assign n15384_o = r[242];
  /* fpu.vhdl:1421:47  */
  assign n15385_o = ~n15384_o;
  /* fpu.vhdl:1421:25  */
  assign n15388_o = n15385_o ? 7'b0101100 : 7'b1001011;
  /* fpu.vhdl:1419:25  */
  assign n15389_o = n15382_o ? 7'b1001010 : n15388_o;
  /* fpu.vhdl:1416:25  */
  assign n15390_o = n15379_o ? n13151_o : n15389_o;
  assign n15391_o = r[136];
  /* fpu.vhdl:1416:25  */
  assign n15392_o = n15379_o ? 1'b1 : n15391_o;
  /* fpu.vhdl:1416:25  */
  assign n15395_o = n15379_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1414:21  */
  assign n15397_o = n15375_o == 2'b01;
  /* fpu.vhdl:1426:21  */
  assign n15400_o = n15375_o == 2'b11;
  /* fpu.vhdl:1429:30  */
  assign n15401_o = r[318:239];
  /* fpu.vhdl:1429:32  */
  assign n15402_o = n15401_o[2];
  assign n15405_o = r[136];
  /* fpu.vhdl:1429:25  */
  assign n15406_o = n15402_o ? 1'b1 : n15405_o;
  /* fpu.vhdl:1429:25  */
  assign n15407_o = n15402_o ? n15367_o : 2'b00;
  /* fpu.vhdl:1429:25  */
  assign n15410_o = n15402_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1428:21  */
  assign n15412_o = n15375_o == 2'b10;
  /* fpu.vhdl:1436:21  */
  assign n15415_o = n15375_o == 2'b00;
  assign n15416_o = {n15415_o, n15412_o, n15400_o, n15397_o};
  /* fpu.vhdl:1413:17  */
  always @*
    case (n15416_o)
      4'b1000: n15418_o = n13151_o;
      4'b0100: n15418_o = n13151_o;
      4'b0010: n15418_o = 7'b1001110;
      4'b0001: n15418_o = n15390_o;
      default: n15418_o = 7'bX;
    endcase
  assign n15419_o = r[136];
  /* fpu.vhdl:1413:17  */
  always @*
    case (n15416_o)
      4'b1000: n15421_o = n15419_o;
      4'b0100: n15421_o = n15406_o;
      4'b0010: n15421_o = n15419_o;
      4'b0001: n15421_o = n15392_o;
      default: n15421_o = 1'bX;
    endcase
  /* fpu.vhdl:1413:17  */
  always @*
    case (n15416_o)
      4'b1000: n15423_o = 2'b10;
      4'b0100: n15423_o = n15407_o;
      4'b0010: n15423_o = n15367_o;
      4'b0001: n15423_o = n15367_o;
      default: n15423_o = 2'bX;
    endcase
  assign n15424_o = r[663:651];
  /* fpu.vhdl:1413:17  */
  always @*
    case (n15416_o)
      4'b1000: n15426_o = n15424_o;
      4'b0100: n15426_o = n15424_o;
      4'b0010: n15426_o = n15424_o;
      4'b0001: n15426_o = n15377_o;
      default: n15426_o = 13'bX;
    endcase
  /* fpu.vhdl:1413:17  */
  always @*
    case (n15416_o)
      4'b1000: n15431_o = 1'b1;
      4'b0100: n15431_o = 1'b1;
      4'b0010: n15431_o = 1'b0;
      4'b0001: n15431_o = 1'b0;
      default: n15431_o = 1'bX;
    endcase
  /* fpu.vhdl:1413:17  */
  always @*
    case (n15416_o)
      4'b1000: n15435_o = 1'b1;
      4'b0100: n15435_o = 1'b0;
      4'b0010: n15435_o = 1'b0;
      4'b0001: n15435_o = 1'b0;
      default: n15435_o = 1'bX;
    endcase
  /* fpu.vhdl:1413:17  */
  always @*
    case (n15416_o)
      4'b1000: n15438_o = 1'b0;
      4'b0100: n15438_o = n15410_o;
      4'b0010: n15438_o = 1'b0;
      4'b0001: n15438_o = n15395_o;
      default: n15438_o = 1'bX;
    endcase
  /* fpu.vhdl:1405:13  */
  assign n15440_o = n13567_o == 7'b0010101;
  /* fpu.vhdl:1446:36  */
  assign n15441_o = r[238:159];
  /* fpu.vhdl:1446:38  */
  assign n15442_o = n15441_o[2];
  /* fpu.vhdl:1447:37  */
  assign n15443_o = r[238:159];
  /* fpu.vhdl:1447:39  */
  assign n15444_o = n15443_o[1:0];
  /* fpu.vhdl:1448:35  */
  assign n15445_o = r[238:159];
  /* fpu.vhdl:1448:37  */
  assign n15446_o = n15445_o[15:3];
  /* fpu.vhdl:1454:29  */
  assign n15452_o = r[238:159];
  /* fpu.vhdl:1454:31  */
  assign n15453_o = n15452_o[2];
  /* fpu.vhdl:1454:46  */
  assign n15454_o = r[398:319];
  /* fpu.vhdl:1454:48  */
  assign n15455_o = n15454_o[2];
  /* fpu.vhdl:1454:40  */
  assign n15456_o = n15453_o ^ n15455_o;
  /* fpu.vhdl:1454:63  */
  assign n15457_o = r[318:239];
  /* fpu.vhdl:1454:65  */
  assign n15458_o = n15457_o[2];
  /* fpu.vhdl:1454:57  */
  assign n15459_o = n15456_o ^ n15458_o;
  /* fpu.vhdl:1454:84  */
  assign n15460_o = r[18];
  /* fpu.vhdl:1454:74  */
  assign n15461_o = n15459_o ^ n15460_o;
  /* fpu.vhdl:1455:22  */
  assign n15462_o = r[238:159];
  /* fpu.vhdl:1455:24  */
  assign n15463_o = n15462_o[1:0];
  /* fpu.vhdl:1455:30  */
  assign n15465_o = n15463_o == 2'b01;
  /* fpu.vhdl:1455:45  */
  assign n15466_o = r[398:319];
  /* fpu.vhdl:1455:47  */
  assign n15467_o = n15466_o[1:0];
  /* fpu.vhdl:1455:53  */
  assign n15469_o = n15467_o == 2'b01;
  /* fpu.vhdl:1455:39  */
  assign n15470_o = n15465_o & n15469_o;
  /* fpu.vhdl:1456:24  */
  assign n15471_o = r[318:239];
  /* fpu.vhdl:1456:26  */
  assign n15472_o = n15471_o[1:0];
  /* fpu.vhdl:1456:32  */
  assign n15474_o = n15472_o == 2'b01;
  /* fpu.vhdl:1456:46  */
  assign n15475_o = r[318:239];
  /* fpu.vhdl:1456:48  */
  assign n15476_o = n15475_o[1:0];
  /* fpu.vhdl:1456:54  */
  assign n15478_o = n15476_o == 2'b00;
  /* fpu.vhdl:1456:41  */
  assign n15479_o = n15474_o | n15478_o;
  /* fpu.vhdl:1455:62  */
  assign n15480_o = n15470_o & n15479_o;
  /* fpu.vhdl:1457:38  */
  assign n15481_o = ~n15461_o;
  /* fpu.vhdl:1458:33  */
  assign n15482_o = r[238:159];
  /* fpu.vhdl:1458:35  */
  assign n15483_o = n15482_o[15:3];
  /* fpu.vhdl:1458:48  */
  assign n15484_o = r[398:319];
  /* fpu.vhdl:1458:50  */
  assign n15485_o = n15484_o[15:3];
  /* fpu.vhdl:1458:44  */
  assign n15486_o = n15483_o + n15485_o;
  /* fpu.vhdl:1461:36  */
  assign n15487_o = r[229];
  /* fpu.vhdl:1461:41  */
  assign n15488_o = ~n15487_o;
  /* fpu.vhdl:1463:39  */
  assign n15490_o = r[389];
  /* fpu.vhdl:1463:44  */
  assign n15491_o = ~n15490_o;
  /* fpu.vhdl:1465:29  */
  assign n15493_o = r[318:239];
  /* fpu.vhdl:1465:31  */
  assign n15494_o = n15493_o[1:0];
  /* fpu.vhdl:1465:37  */
  assign n15496_o = n15494_o == 2'b00;
  /* fpu.vhdl:1467:44  */
  assign n15497_o = r[238:159];
  /* fpu.vhdl:1467:46  */
  assign n15498_o = n15497_o[2];
  /* fpu.vhdl:1467:61  */
  assign n15499_o = r[398:319];
  /* fpu.vhdl:1467:63  */
  assign n15500_o = n15499_o[2];
  /* fpu.vhdl:1467:55  */
  assign n15501_o = n15498_o ^ n15500_o;
  /* fpu.vhdl:1467:82  */
  assign n15502_o = r[19];
  /* fpu.vhdl:1467:72  */
  assign n15503_o = n15501_o ^ n15502_o;
  /* fpu.vhdl:1471:29  */
  assign n15507_o = r[705];
  /* fpu.vhdl:1471:38  */
  assign n15508_o = ~n15507_o;
  /* fpu.vhdl:1473:49  */
  assign n15509_o = r[318:239];
  /* fpu.vhdl:1473:51  */
  assign n15510_o = n15509_o[2];
  /* fpu.vhdl:1473:70  */
  assign n15511_o = r[18];
  /* fpu.vhdl:1473:60  */
  assign n15512_o = n15510_o ^ n15511_o;
  /* fpu.vhdl:1473:84  */
  assign n15513_o = r[19];
  /* fpu.vhdl:1473:74  */
  assign n15514_o = n15512_o ^ n15513_o;
  /* fpu.vhdl:1473:42  */
  assign n15515_o = ~n15514_o;
  /* fpu.vhdl:1479:38  */
  assign n15518_o = r[318:239];
  /* fpu.vhdl:1479:40  */
  assign n15519_o = n15518_o[15:3];
  /* fpu.vhdl:1479:49  */
  assign n15520_o = n15519_o - n15486_o;
  /* fpu.vhdl:1479:58  */
  assign n15522_o = n15520_o + 13'b0000001000000;
  /* fpu.vhdl:1481:49  */
  assign n15523_o = r[238:159];
  /* fpu.vhdl:1481:51  */
  assign n15524_o = n15523_o[2];
  /* fpu.vhdl:1481:66  */
  assign n15525_o = r[398:319];
  /* fpu.vhdl:1481:68  */
  assign n15526_o = n15525_o[2];
  /* fpu.vhdl:1481:60  */
  assign n15527_o = n15524_o ^ n15526_o;
  /* fpu.vhdl:1481:87  */
  assign n15528_o = r[19];
  /* fpu.vhdl:1481:77  */
  assign n15529_o = n15527_o ^ n15528_o;
  /* fpu.vhdl:1481:91  */
  assign n15530_o = n15529_o ^ n15461_o;
  /* fpu.vhdl:1481:42  */
  assign n15531_o = ~n15530_o;
  /* fpu.vhdl:1482:43  */
  assign n15532_o = r[318:239];
  /* fpu.vhdl:1482:45  */
  assign n15533_o = n15532_o[15:3];
  /* fpu.vhdl:1471:21  */
  assign n15535_o = n15508_o ? 1'b1 : 1'b0;
  assign n15536_o = {n15522_o, n15533_o};
  /* fpu.vhdl:1471:21  */
  assign n15537_o = n15508_o ? 7'b0011111 : 7'b0100000;
  /* fpu.vhdl:1471:21  */
  assign n15538_o = n15508_o ? n15515_o : n15531_o;
  assign n15539_o = {13'b0000000000000, n15486_o};
  /* fpu.vhdl:1471:21  */
  assign n15540_o = n15508_o ? n15539_o : n15536_o;
  /* fpu.vhdl:1465:21  */
  assign n15541_o = n15496_o ? 1'b1 : n15535_o;
  /* fpu.vhdl:1465:21  */
  assign n15542_o = n15496_o ? 7'b0011110 : n15537_o;
  /* fpu.vhdl:1465:21  */
  assign n15543_o = n15496_o ? n15503_o : n15538_o;
  assign n15544_o = {13'b0000000000000, n15486_o};
  /* fpu.vhdl:1465:21  */
  assign n15545_o = n15496_o ? n15544_o : n15540_o;
  assign n15546_o = n13465_o[10];
  assign n15547_o = r[707];
  /* fpu.vhdl:650:9  */
  assign n15548_o = n13152_o ? n15546_o : n15547_o;
  /* fpu.vhdl:1465:21  */
  assign n15549_o = n15496_o ? 1'b1 : n15548_o;
  /* fpu.vhdl:1463:21  */
  assign n15550_o = n15491_o ? 1'b0 : n15541_o;
  /* fpu.vhdl:1463:21  */
  assign n15551_o = n15491_o ? 7'b1001100 : n15542_o;
  /* fpu.vhdl:1463:21  */
  assign n15552_o = n15491_o ? n15442_o : n15543_o;
  assign n15553_o = {13'b0000000000000, n15486_o};
  /* fpu.vhdl:1463:21  */
  assign n15554_o = n15491_o ? n15553_o : n15545_o;
  assign n15555_o = n13465_o[10];
  assign n15556_o = r[707];
  /* fpu.vhdl:650:9  */
  assign n15557_o = n13152_o ? n15555_o : n15556_o;
  /* fpu.vhdl:1463:21  */
  assign n15558_o = n15491_o ? n15557_o : n15549_o;
  /* fpu.vhdl:1461:21  */
  assign n15559_o = n15488_o ? 1'b0 : n15550_o;
  /* fpu.vhdl:1461:21  */
  assign n15560_o = n15488_o ? 7'b1001000 : n15551_o;
  /* fpu.vhdl:1461:21  */
  assign n15561_o = n15488_o ? n15442_o : n15552_o;
  assign n15562_o = {13'b0000000000000, n15486_o};
  /* fpu.vhdl:1461:21  */
  assign n15563_o = n15488_o ? n15562_o : n15554_o;
  assign n15564_o = n13465_o[10];
  assign n15565_o = r[707];
  /* fpu.vhdl:650:9  */
  assign n15566_o = n13152_o ? n15564_o : n15565_o;
  /* fpu.vhdl:1461:21  */
  assign n15567_o = n15488_o ? n15566_o : n15558_o;
  /* fpu.vhdl:1486:26  */
  assign n15568_o = r[238:159];
  /* fpu.vhdl:1486:28  */
  assign n15569_o = n15568_o[1:0];
  /* fpu.vhdl:1486:34  */
  assign n15571_o = n15569_o == 2'b11;
  /* fpu.vhdl:1486:45  */
  assign n15572_o = r[318:239];
  /* fpu.vhdl:1486:47  */
  assign n15573_o = n15572_o[1:0];
  /* fpu.vhdl:1486:53  */
  assign n15575_o = n15573_o == 2'b11;
  /* fpu.vhdl:1486:40  */
  assign n15576_o = n15571_o | n15575_o;
  /* fpu.vhdl:1486:64  */
  assign n15577_o = r[398:319];
  /* fpu.vhdl:1486:66  */
  assign n15578_o = n15577_o[1:0];
  /* fpu.vhdl:1486:72  */
  assign n15580_o = n15578_o == 2'b11;
  /* fpu.vhdl:1486:59  */
  assign n15581_o = n15576_o | n15580_o;
  /* fpu.vhdl:1488:30  */
  assign n15583_o = r[238:159];
  /* fpu.vhdl:1488:32  */
  assign n15584_o = n15583_o[1:0];
  /* fpu.vhdl:1488:38  */
  assign n15586_o = n15584_o == 2'b00;
  /* fpu.vhdl:1488:51  */
  assign n15587_o = r[398:319];
  /* fpu.vhdl:1488:53  */
  assign n15588_o = n15587_o[1:0];
  /* fpu.vhdl:1488:59  */
  assign n15590_o = n15588_o == 2'b10;
  /* fpu.vhdl:1488:45  */
  assign n15591_o = n15586_o & n15590_o;
  /* fpu.vhdl:1489:28  */
  assign n15592_o = r[238:159];
  /* fpu.vhdl:1489:30  */
  assign n15593_o = n15592_o[1:0];
  /* fpu.vhdl:1489:36  */
  assign n15595_o = n15593_o == 2'b10;
  /* fpu.vhdl:1489:53  */
  assign n15596_o = r[398:319];
  /* fpu.vhdl:1489:55  */
  assign n15597_o = n15596_o[1:0];
  /* fpu.vhdl:1489:61  */
  assign n15599_o = n15597_o == 2'b00;
  /* fpu.vhdl:1489:47  */
  assign n15600_o = n15595_o & n15599_o;
  /* fpu.vhdl:1488:71  */
  assign n15601_o = n15591_o | n15600_o;
  /* fpu.vhdl:1493:29  */
  assign n15603_o = r[238:159];
  /* fpu.vhdl:1493:31  */
  assign n15604_o = n15603_o[1:0];
  /* fpu.vhdl:1493:37  */
  assign n15606_o = n15604_o == 2'b10;
  /* fpu.vhdl:1493:53  */
  assign n15607_o = r[398:319];
  /* fpu.vhdl:1493:55  */
  assign n15608_o = n15607_o[1:0];
  /* fpu.vhdl:1493:61  */
  assign n15610_o = n15608_o == 2'b10;
  /* fpu.vhdl:1493:48  */
  assign n15611_o = n15606_o | n15610_o;
  /* fpu.vhdl:1494:30  */
  assign n15612_o = r[318:239];
  /* fpu.vhdl:1494:32  */
  assign n15613_o = n15612_o[1:0];
  /* fpu.vhdl:1494:38  */
  assign n15615_o = n15613_o == 2'b10;
  /* fpu.vhdl:1494:60  */
  assign n15616_o = ~n15461_o;
  /* fpu.vhdl:1494:49  */
  assign n15617_o = n15615_o & n15616_o;
  /* fpu.vhdl:1501:48  */
  assign n15620_o = r[238:159];
  /* fpu.vhdl:1501:50  */
  assign n15621_o = n15620_o[2];
  /* fpu.vhdl:1501:65  */
  assign n15622_o = r[398:319];
  /* fpu.vhdl:1501:67  */
  assign n15623_o = n15622_o[2];
  /* fpu.vhdl:1501:59  */
  assign n15624_o = n15621_o ^ n15623_o;
  /* fpu.vhdl:1501:86  */
  assign n15625_o = r[19];
  /* fpu.vhdl:1501:76  */
  assign n15626_o = n15624_o ^ n15625_o;
  assign n15627_o = {2'b10, n15626_o};
  assign n15628_o = r[150];
  /* fpu.vhdl:1493:21  */
  assign n15629_o = n15660_o ? 1'b1 : n15628_o;
  assign n15630_o = {n15444_o, n15442_o};
  /* fpu.vhdl:1494:25  */
  assign n15631_o = n15617_o ? n15630_o : n15627_o;
  /* fpu.vhdl:1494:25  */
  assign n15634_o = n15617_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:1494:25  */
  assign n15637_o = n15617_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1508:30  */
  assign n15639_o = r[318:239];
  /* fpu.vhdl:1508:32  */
  assign n15640_o = n15639_o[1:0];
  /* fpu.vhdl:1508:38  */
  assign n15642_o = n15640_o != 2'b00;
  /* fpu.vhdl:1508:46  */
  assign n15643_o = n15642_o | n15461_o;
  /* fpu.vhdl:1509:52  */
  assign n15644_o = r[18];
  /* fpu.vhdl:1509:66  */
  assign n15645_o = r[19];
  /* fpu.vhdl:1509:56  */
  assign n15646_o = n15644_o ^ n15645_o;
  /* fpu.vhdl:1509:41  */
  assign n15647_o = ~n15646_o;
  /* fpu.vhdl:1512:43  */
  assign n15648_o = r[318:239];
  /* fpu.vhdl:1512:45  */
  assign n15649_o = n15648_o[2];
  /* fpu.vhdl:1512:71  */
  assign n15650_o = r[701];
  /* fpu.vhdl:1512:91  */
  assign n15651_o = r[700];
  /* fpu.vhdl:1512:75  */
  assign n15652_o = n15650_o & n15651_o;
  /* fpu.vhdl:1512:54  */
  assign n15653_o = n15649_o ^ n15652_o;
  /* fpu.vhdl:1512:106  */
  assign n15654_o = r[19];
  /* fpu.vhdl:1512:96  */
  assign n15655_o = n15653_o ^ n15654_o;
  /* fpu.vhdl:1508:25  */
  assign n15656_o = n15643_o ? n15647_o : n15655_o;
  /* fpu.vhdl:1493:21  */
  assign n15658_o = n15611_o ? n13151_o : 7'b1001111;
  /* fpu.vhdl:1493:21  */
  assign n15660_o = n15611_o & n15617_o;
  assign n15661_o = {n15444_o, n15442_o};
  /* fpu.vhdl:1493:21  */
  assign n15662_o = n15611_o ? n15631_o : n15661_o;
  /* fpu.vhdl:1493:21  */
  assign n15663_o = n15611_o ? 2'b00 : 2'b10;
  assign n15664_o = r[720];
  /* fpu.vhdl:1493:21  */
  assign n15665_o = n15611_o ? n15664_o : n15656_o;
  /* fpu.vhdl:1493:21  */
  assign n15667_o = n15611_o ? n15634_o : 1'b0;
  /* fpu.vhdl:1493:21  */
  assign n15669_o = n15611_o ? n15637_o : 1'b0;
  /* fpu.vhdl:1488:21  */
  assign n15670_o = n15601_o ? n13151_o : n15658_o;
  assign n15671_o = r[147];
  /* fpu.vhdl:1488:21  */
  assign n15672_o = n15601_o ? 1'b1 : n15671_o;
  assign n15673_o = r[150];
  /* fpu.vhdl:1488:21  */
  assign n15674_o = n15601_o ? n15673_o : n15629_o;
  assign n15675_o = {n15444_o, n15442_o};
  /* fpu.vhdl:1488:21  */
  assign n15676_o = n15601_o ? n15675_o : n15662_o;
  /* fpu.vhdl:1488:21  */
  assign n15677_o = n15601_o ? 2'b00 : n15663_o;
  assign n15678_o = r[720];
  /* fpu.vhdl:1488:21  */
  assign n15679_o = n15601_o ? n15678_o : n15665_o;
  /* fpu.vhdl:1488:21  */
  assign n15681_o = n15601_o ? 1'b0 : n15667_o;
  /* fpu.vhdl:1488:21  */
  assign n15683_o = n15601_o ? 1'b1 : n15669_o;
  /* fpu.vhdl:1486:21  */
  assign n15684_o = n15581_o ? 7'b1001110 : n15670_o;
  assign n15685_o = r[147];
  /* fpu.vhdl:1486:21  */
  assign n15686_o = n15581_o ? n15685_o : n15672_o;
  assign n15687_o = r[150];
  /* fpu.vhdl:1486:21  */
  assign n15688_o = n15581_o ? n15687_o : n15674_o;
  assign n15689_o = {n15444_o, n15442_o};
  /* fpu.vhdl:1486:21  */
  assign n15690_o = n15581_o ? n15689_o : n15676_o;
  /* fpu.vhdl:1486:21  */
  assign n15691_o = n15581_o ? 2'b00 : n15677_o;
  assign n15692_o = r[720];
  /* fpu.vhdl:1486:21  */
  assign n15693_o = n15581_o ? n15692_o : n15679_o;
  /* fpu.vhdl:1486:21  */
  assign n15695_o = n15581_o ? 1'b0 : n15681_o;
  /* fpu.vhdl:1486:21  */
  assign n15697_o = n15581_o ? 1'b0 : n15683_o;
  /* fpu.vhdl:1455:17  */
  assign n15698_o = n15480_o ? n15559_o : 1'b0;
  /* fpu.vhdl:1455:17  */
  assign n15699_o = n15480_o ? n15560_o : n15684_o;
  assign n15700_o = r[147];
  /* fpu.vhdl:1455:17  */
  assign n15701_o = n15480_o ? n15700_o : n15686_o;
  assign n15702_o = r[150];
  /* fpu.vhdl:1455:17  */
  assign n15703_o = n15480_o ? n15702_o : n15688_o;
  assign n15704_o = n15690_o[0];
  /* fpu.vhdl:1455:17  */
  assign n15705_o = n15480_o ? n15561_o : n15704_o;
  assign n15706_o = n15690_o[2:1];
  /* fpu.vhdl:1455:17  */
  assign n15707_o = n15480_o ? n15444_o : n15706_o;
  assign n15708_o = {13'b0000000000000, n15446_o};
  /* fpu.vhdl:1455:17  */
  assign n15709_o = n15480_o ? n15563_o : n15708_o;
  assign n15710_o = n13465_o[6];
  assign n15711_o = r[703];
  /* fpu.vhdl:650:9  */
  assign n15712_o = n13152_o ? n15710_o : n15711_o;
  /* fpu.vhdl:1455:17  */
  assign n15713_o = n15480_o ? n15481_o : n15712_o;
  assign n15714_o = n13465_o[10];
  assign n15715_o = r[707];
  /* fpu.vhdl:650:9  */
  assign n15716_o = n13152_o ? n15714_o : n15715_o;
  /* fpu.vhdl:1455:17  */
  assign n15717_o = n15480_o ? n15567_o : n15716_o;
  /* fpu.vhdl:1455:17  */
  assign n15718_o = n15480_o ? 2'b00 : n15691_o;
  assign n15719_o = r[720];
  /* fpu.vhdl:1455:17  */
  assign n15720_o = n15480_o ? n15719_o : n15693_o;
  /* fpu.vhdl:1455:17  */
  assign n15722_o = n15480_o ? 1'b0 : n15695_o;
  /* fpu.vhdl:1455:17  */
  assign n15724_o = n15480_o ? 1'b0 : n15697_o;
  /* fpu.vhdl:1442:13  */
  assign n15727_o = n13567_o == 7'b0010011;
  /* fpu.vhdl:1521:26  */
  assign n15729_o = r[21];
  /* fpu.vhdl:1521:17  */
  assign n15732_o = n15729_o ? 2'b11 : 2'b10;
  /* fpu.vhdl:1518:13  */
  assign n15734_o = n13567_o == 7'b1001000;
  /* fpu.vhdl:1531:26  */
  assign n15735_o = r[21];
  /* fpu.vhdl:1532:36  */
  assign n15736_o = r[389];
  /* fpu.vhdl:1533:34  */
  assign n15737_o = r[20];
  /* fpu.vhdl:1533:38  */
  assign n15738_o = ~n15737_o;
  /* fpu.vhdl:1533:49  */
  assign n15739_o = r[318:239];
  /* fpu.vhdl:1533:51  */
  assign n15740_o = n15739_o[1:0];
  /* fpu.vhdl:1533:57  */
  assign n15742_o = n15740_o == 2'b00;
  /* fpu.vhdl:1533:44  */
  assign n15743_o = n15738_o | n15742_o;
  /* fpu.vhdl:1538:40  */
  assign n15748_o = n13526_o + 13'b0000000000001;
  /* fpu.vhdl:1538:49  */
  assign n15749_o = r[318:239];
  /* fpu.vhdl:1538:51  */
  assign n15750_o = n15749_o[15:3];
  /* fpu.vhdl:1538:44  */
  assign n15751_o = $signed(n15748_o) >= $signed(n15750_o);
  /* fpu.vhdl:1538:29  */
  assign n15753_o = n15751_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1533:25  */
  assign n15756_o = n15743_o ? 7'b0011110 : 7'b0010011;
  assign n15757_o = n13465_o[8];
  assign n15758_o = r[705];
  /* fpu.vhdl:650:9  */
  assign n15759_o = n13152_o ? n15757_o : n15758_o;
  /* fpu.vhdl:1533:25  */
  assign n15760_o = n15743_o ? n15759_o : n15753_o;
  /* fpu.vhdl:1532:21  */
  assign n15761_o = n15769_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1533:25  */
  assign n15762_o = n15743_o ? 2'b00 : 2'b10;
  /* fpu.vhdl:1532:21  */
  assign n15764_o = n15736_o ? n15756_o : 7'b1001100;
  assign n15765_o = n13465_o[8];
  assign n15766_o = r[705];
  /* fpu.vhdl:650:9  */
  assign n15767_o = n13152_o ? n15765_o : n15766_o;
  /* fpu.vhdl:1532:21  */
  assign n15768_o = n15736_o ? n15760_o : n15767_o;
  /* fpu.vhdl:1532:21  */
  assign n15769_o = n15736_o & n15743_o;
  /* fpu.vhdl:1531:17  */
  assign n15770_o = n15783_o ? n15762_o : 2'b00;
  /* fpu.vhdl:1548:36  */
  assign n15771_o = r[309];
  /* fpu.vhdl:1548:21  */
  assign n15775_o = n15771_o ? 7'b0100110 : 7'b1001010;
  /* fpu.vhdl:1548:21  */
  assign n15776_o = n15771_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1531:17  */
  assign n15777_o = n15735_o ? n15764_o : n15775_o;
  assign n15778_o = n13465_o[8];
  assign n15779_o = r[705];
  /* fpu.vhdl:650:9  */
  assign n15780_o = n13152_o ? n15778_o : n15779_o;
  /* fpu.vhdl:1531:17  */
  assign n15781_o = n15735_o ? n15768_o : n15780_o;
  /* fpu.vhdl:1531:17  */
  assign n15782_o = n15735_o ? n15761_o : n15776_o;
  /* fpu.vhdl:1531:17  */
  assign n15783_o = n15735_o & n15736_o;
  /* fpu.vhdl:1527:13  */
  assign n15785_o = n13567_o == 7'b1001001;
  /* fpu.vhdl:1558:34  */
  assign n15786_o = r[708];
  /* fpu.vhdl:1556:13  */
  assign n15789_o = n13567_o == 7'b1001010;
  /* fpu.vhdl:1563:22  */
  assign n15790_o = r[708];
  /* fpu.vhdl:1563:30  */
  assign n15791_o = ~n15790_o;
  /* fpu.vhdl:1564:39  */
  assign n15792_o = r[663:651];
  /* fpu.vhdl:1564:54  */
  assign n15793_o = r[676:664];
  /* fpu.vhdl:1564:50  */
  assign n15794_o = n15792_o + n15793_o;
  /* fpu.vhdl:1563:17  */
  assign n15795_o = n15791_o ? n15794_o : n13526_o;
  /* fpu.vhdl:1561:13  */
  assign n15799_o = n13567_o == 7'b1001011;
  /* fpu.vhdl:1571:13  */
  assign n15802_o = n13567_o == 7'b1001100;
  /* fpu.vhdl:1578:26  */
  assign n15803_o = r[20];
  /* fpu.vhdl:1578:30  */
  assign n15804_o = ~n15803_o;
  /* fpu.vhdl:1578:41  */
  assign n15805_o = r[318:239];
  /* fpu.vhdl:1578:43  */
  assign n15806_o = n15805_o[1:0];
  /* fpu.vhdl:1578:49  */
  assign n15808_o = n15806_o == 2'b00;
  /* fpu.vhdl:1578:36  */
  assign n15809_o = n15804_o | n15808_o;
  /* fpu.vhdl:1583:32  */
  assign n15814_o = n13526_o + 13'b0000000000001;
  /* fpu.vhdl:1583:41  */
  assign n15815_o = r[318:239];
  /* fpu.vhdl:1583:43  */
  assign n15816_o = n15815_o[15:3];
  /* fpu.vhdl:1583:36  */
  assign n15817_o = $signed(n15814_o) >= $signed(n15816_o);
  /* fpu.vhdl:1583:21  */
  assign n15819_o = n15817_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1578:17  */
  assign n15822_o = n15809_o ? 7'b0011110 : 7'b0010011;
  assign n15823_o = n13465_o[8];
  assign n15824_o = r[705];
  /* fpu.vhdl:650:9  */
  assign n15825_o = n13152_o ? n15823_o : n15824_o;
  /* fpu.vhdl:1578:17  */
  assign n15826_o = n15809_o ? n15825_o : n15819_o;
  /* fpu.vhdl:1578:17  */
  assign n15827_o = n15809_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1578:17  */
  assign n15828_o = n15809_o ? 2'b00 : 2'b10;
  /* fpu.vhdl:1575:13  */
  assign n15830_o = n13567_o == 7'b1001101;
  /* fpu.vhdl:1592:30  */
  assign n15831_o = r[318:239];
  /* fpu.vhdl:1592:32  */
  assign n15832_o = n15831_o[15:3];
  /* fpu.vhdl:1592:45  */
  assign n15833_o = r[238:159];
  /* fpu.vhdl:1592:47  */
  assign n15834_o = n15833_o[15:3];
  /* fpu.vhdl:1592:41  */
  assign n15835_o = n15832_o - n15834_o;
  /* fpu.vhdl:1593:35  */
  assign n15836_o = r[318:239];
  /* fpu.vhdl:1593:37  */
  assign n15837_o = n15836_o[15:3];
  /* fpu.vhdl:1590:13  */
  assign n15841_o = n13567_o == 7'b0011000;
  /* fpu.vhdl:1602:33  */
  assign n15842_o = r[126];
  /* fpu.vhdl:1603:22  */
  assign n15843_o = r[706];
  /* fpu.vhdl:1603:17  */
  assign n15846_o = n15843_o ? 2'b01 : 2'b10;
  /* fpu.vhdl:1597:13  */
  assign n15849_o = n13567_o == 7'b0011001;
  /* fpu.vhdl:1613:33  */
  assign n15850_o = r[703];
  /* fpu.vhdl:1614:31  */
  assign n15851_o = r[703];
  /* fpu.vhdl:1614:53  */
  assign n15852_o = r[519];
  /* fpu.vhdl:1614:47  */
  assign n15853_o = ~n15852_o;
  /* fpu.vhdl:1614:43  */
  assign n15854_o = n15851_o & n15853_o;
  /* fpu.vhdl:1610:13  */
  assign n15858_o = n13567_o == 7'b0011010;
  /* fpu.vhdl:1621:23  */
  assign n15859_o = r[462];
  /* fpu.vhdl:1623:44  */
  assign n15860_o = r[648];
  /* fpu.vhdl:1623:38  */
  assign n15861_o = ~n15860_o;
  /* fpu.vhdl:1627:26  */
  assign n15863_o = r[454];
  /* fpu.vhdl:1631:21  */
  assign n15866_o = n13535_o ? 7'b1000011 : 7'b1000100;
  /* fpu.vhdl:1636:26  */
  assign n15867_o = r[453];
  /* fpu.vhdl:1639:32  */
  assign n15869_o = r_hi_nz | r_lo_nz;
  /* fpu.vhdl:1639:49  */
  assign n15870_o = r[400];
  /* fpu.vhdl:1639:43  */
  assign n15871_o = n15869_o | n15870_o;
  /* fpu.vhdl:1639:59  */
  assign n15872_o = r[399];
  /* fpu.vhdl:1639:53  */
  assign n15873_o = n15871_o | n15872_o;
  /* fpu.vhdl:1639:64  */
  assign n15874_o = ~n15873_o;
  /* fpu.vhdl:1642:26  */
  assign n15876_o = r[703];
  /* fpu.vhdl:1644:54  */
  assign n15877_o = r[701];
  /* fpu.vhdl:1644:74  */
  assign n15878_o = r[700];
  /* fpu.vhdl:1644:58  */
  assign n15879_o = n15877_o & n15878_o;
  assign n15880_o = r[648];
  /* fpu.vhdl:1642:21  */
  assign n15881_o = n15876_o ? n15879_o : n15880_o;
  assign n15883_o = {2'b00, n15881_o};
  /* fpu.vhdl:1639:17  */
  assign n15884_o = n15874_o ? n13151_o : 7'b1000001;
  assign n15885_o = r[650:648];
  /* fpu.vhdl:1639:17  */
  assign n15886_o = n15874_o ? n15883_o : n15885_o;
  /* fpu.vhdl:1639:17  */
  assign n15889_o = n15874_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1639:17  */
  assign n15892_o = n15874_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:1636:17  */
  assign n15893_o = n15867_o ? 7'b1000100 : n15884_o;
  assign n15894_o = r[650:648];
  /* fpu.vhdl:1636:17  */
  assign n15895_o = n15867_o ? n15894_o : n15886_o;
  /* fpu.vhdl:1636:17  */
  assign n15897_o = n15867_o ? 1'b0 : n15889_o;
  /* fpu.vhdl:1636:17  */
  assign n15899_o = n15867_o ? 1'b0 : n15892_o;
  /* fpu.vhdl:1636:17  */
  assign n15902_o = n15867_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1627:17  */
  assign n15905_o = n15863_o ? 2'b01 : 2'b00;
  /* fpu.vhdl:1627:17  */
  assign n15906_o = n15863_o ? n15866_o : n15893_o;
  assign n15907_o = r[650:648];
  /* fpu.vhdl:1627:17  */
  assign n15908_o = n15863_o ? n15907_o : n15895_o;
  /* fpu.vhdl:1627:17  */
  assign n15910_o = n15863_o ? 1'b0 : n15897_o;
  /* fpu.vhdl:1627:17  */
  assign n15912_o = n15863_o ? 1'b0 : n15899_o;
  /* fpu.vhdl:1627:17  */
  assign n15914_o = n15863_o ? 1'b1 : n15902_o;
  /* fpu.vhdl:1621:17  */
  assign n15916_o = n15859_o ? 2'b00 : n15905_o;
  /* fpu.vhdl:1621:17  */
  assign n15919_o = n15859_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1621:17  */
  assign n15922_o = n15859_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1621:17  */
  assign n15923_o = n15859_o ? 7'b1000000 : n15906_o;
  assign n15924_o = n15908_o[0];
  /* fpu.vhdl:1621:17  */
  assign n15925_o = n15859_o ? n15861_o : n15924_o;
  assign n15926_o = n15908_o[2:1];
  assign n15927_o = r[650:649];
  /* fpu.vhdl:1621:17  */
  assign n15928_o = n15859_o ? n15927_o : n15926_o;
  /* fpu.vhdl:1621:17  */
  assign n15930_o = n15859_o ? 1'b0 : n15910_o;
  /* fpu.vhdl:1621:17  */
  assign n15932_o = n15859_o ? 1'b0 : n15912_o;
  /* fpu.vhdl:1621:17  */
  assign n15934_o = n15859_o ? 1'b0 : n15914_o;
  /* fpu.vhdl:1618:13  */
  assign n15936_o = n13567_o == 7'b0011011;
  /* fpu.vhdl:1652:13  */
  assign n15939_o = n13567_o == 7'b0011100;
  /* fpu.vhdl:1660:23  */
  assign n15940_o = r[462];
  /* fpu.vhdl:1662:42  */
  assign n15941_o = r[238:159];
  /* fpu.vhdl:1662:44  */
  assign n15942_o = n15941_o[2];
  /* fpu.vhdl:1662:36  */
  assign n15943_o = ~n15942_o;
  /* fpu.vhdl:1662:57  */
  assign n15944_o = r[238:159];
  /* fpu.vhdl:1662:59  */
  assign n15945_o = n15944_o[2];
  /* fpu.vhdl:1662:53  */
  assign n15946_o = {n15943_o, n15945_o};
  /* fpu.vhdl:1662:68  */
  assign n15948_o = {n15946_o, 2'b00};
  /* fpu.vhdl:1663:32  */
  assign n15949_o = r_hi_nz | r_lo_nz;
  /* fpu.vhdl:1663:44  */
  assign n15950_o = ~n15949_o;
  /* fpu.vhdl:1666:38  */
  assign n15952_o = r[238:159];
  /* fpu.vhdl:1666:40  */
  assign n15953_o = n15952_o[2];
  /* fpu.vhdl:1666:57  */
  assign n15954_o = r[238:159];
  /* fpu.vhdl:1666:59  */
  assign n15955_o = n15954_o[2];
  /* fpu.vhdl:1666:51  */
  assign n15956_o = ~n15955_o;
  /* fpu.vhdl:1666:49  */
  assign n15957_o = {n15953_o, n15956_o};
  /* fpu.vhdl:1666:68  */
  assign n15959_o = {n15957_o, 2'b00};
  /* fpu.vhdl:1663:17  */
  assign n15960_o = n15950_o ? 4'b0010 : n15959_o;
  /* fpu.vhdl:1660:17  */
  assign n15961_o = n15940_o ? n15948_o : n15960_o;
  assign n15962_o = {n13479_o, n13564_o, 2'b00, n13477_o, n13562_o, 1'b0, n13475_o, 1'b0, n13558_o, n13473_o, n15961_o, n13471_o, 1'b0, 13'b0000000000000, n13560_o, n13469_o, n13483_o, n13467_o, n13556_o, 1'b0, 1'b0, n13151_o};
  /* fpu.vhdl:1668:56  */
  assign n15963_o = n15962_o[682:679];
  /* fpu.vhdl:1659:13  */
  assign n15967_o = n13567_o == 7'b0011101;
  /* fpu.vhdl:1673:42  */
  assign n15968_o = r[709];
  /* fpu.vhdl:1675:34  */
  assign n15969_o = multiply_to_f[0];
  /* fpu.vhdl:1675:17  */
  assign n15971_o = n15969_o ? 7'b1000000 : n13151_o;
  /* fpu.vhdl:1672:13  */
  assign n15973_o = n13567_o == 7'b0011110;
  /* fpu.vhdl:1681:41  */
  assign n15974_o = r[318:239];
  /* fpu.vhdl:1681:43  */
  assign n15975_o = n15974_o[2];
  /* fpu.vhdl:1681:62  */
  assign n15976_o = r[18];
  /* fpu.vhdl:1681:52  */
  assign n15977_o = n15975_o ^ n15976_o;
  /* fpu.vhdl:1681:76  */
  assign n15978_o = r[19];
  /* fpu.vhdl:1681:66  */
  assign n15979_o = n15977_o ^ n15978_o;
  /* fpu.vhdl:1681:34  */
  assign n15980_o = ~n15979_o;
  /* fpu.vhdl:1683:30  */
  assign n15981_o = r[663:651];
  /* fpu.vhdl:1683:45  */
  assign n15982_o = r[318:239];
  /* fpu.vhdl:1683:47  */
  assign n15983_o = n15982_o[15:3];
  /* fpu.vhdl:1683:41  */
  assign n15984_o = n15981_o - n15983_o;
  /* fpu.vhdl:1687:42  */
  assign n15985_o = r[709];
  /* fpu.vhdl:1688:34  */
  assign n15986_o = multiply_to_f[0];
  /* fpu.vhdl:1688:17  */
  assign n15989_o = n15986_o ? 7'b0011001 : n13151_o;
  /* fpu.vhdl:1688:17  */
  assign n15990_o = n15986_o ? 1'b0 : n13479_o;
  /* fpu.vhdl:1679:13  */
  assign n15992_o = n13567_o == 7'b0011111;
  /* fpu.vhdl:1698:30  */
  assign n15993_o = r[676:664];
  /* fpu.vhdl:1698:36  */
  assign n15995_o = n15993_o - 13'b0000001000000;
  /* fpu.vhdl:1693:13  */
  assign n15998_o = n13567_o == 7'b0100000;
  /* fpu.vhdl:1701:13  */
  assign n16002_o = n13567_o == 7'b0100001;
  /* fpu.vhdl:1709:42  */
  assign n16003_o = r[709];
  /* fpu.vhdl:1710:31  */
  assign n16004_o = r[703];
  /* fpu.vhdl:1714:34  */
  assign n16005_o = multiply_to_f[0];
  /* fpu.vhdl:1714:17  */
  assign n16007_o = n16005_o ? 7'b0100011 : n13151_o;
  /* fpu.vhdl:1707:13  */
  assign n16009_o = n13567_o == 7'b0100010;
  /* fpu.vhdl:1720:23  */
  assign n16010_o = r[462];
  /* fpu.vhdl:1721:44  */
  assign n16011_o = r[648];
  /* fpu.vhdl:1721:38  */
  assign n16012_o = ~n16011_o;
  /* fpu.vhdl:1723:48  */
  assign n16013_o = r[519];
  /* fpu.vhdl:1723:43  */
  assign n16014_o = s_nz | n16013_o;
  /* fpu.vhdl:1723:33  */
  assign n16015_o = ~n16014_o;
  /* fpu.vhdl:1720:17  */
  assign n16018_o = n16010_o ? 2'b01 : 2'b00;
  /* fpu.vhdl:1720:17  */
  assign n16021_o = n16010_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1720:17  */
  assign n16023_o = n16010_o ? n16015_o : 1'b0;
  assign n16024_o = r[648];
  /* fpu.vhdl:1720:17  */
  assign n16025_o = n16010_o ? n16012_o : n16024_o;
  /* fpu.vhdl:1720:17  */
  assign n16028_o = n16010_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1718:13  */
  assign n16032_o = n13567_o == 7'b0100011;
  /* fpu.vhdl:1732:24  */
  assign n16033_o = r[455];
  /* fpu.vhdl:1732:29  */
  assign n16034_o = n16033_o | r_hi_nz;
  /* fpu.vhdl:1732:40  */
  assign n16035_o = n16034_o | r_lo_nz;
  /* fpu.vhdl:1732:57  */
  assign n16036_o = r[400];
  /* fpu.vhdl:1732:51  */
  assign n16037_o = n16035_o | n16036_o;
  /* fpu.vhdl:1732:67  */
  assign n16038_o = r[399];
  /* fpu.vhdl:1732:61  */
  assign n16039_o = n16037_o | n16038_o;
  /* fpu.vhdl:1732:72  */
  assign n16040_o = ~n16039_o;
  /* fpu.vhdl:1733:29  */
  assign n16041_o = ~s_nz;
  /* fpu.vhdl:1736:54  */
  assign n16043_o = r[701];
  /* fpu.vhdl:1736:74  */
  assign n16044_o = r[700];
  /* fpu.vhdl:1736:58  */
  assign n16045_o = n16043_o & n16044_o;
  /* fpu.vhdl:1733:21  */
  assign n16048_o = n16041_o ? 2'b00 : 2'b01;
  assign n16049_o = {2'b00, n16045_o};
  assign n16050_o = r[650:648];
  /* fpu.vhdl:1732:17  */
  assign n16051_o = n16071_o ? n16049_o : n16050_o;
  /* fpu.vhdl:1733:21  */
  assign n16054_o = n16041_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1733:21  */
  assign n16057_o = n16041_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:1745:26  */
  assign n16058_o = r[455:453];
  /* fpu.vhdl:1745:41  */
  assign n16060_o = n16058_o == 3'b001;
  /* fpu.vhdl:1745:17  */
  assign n16063_o = n16060_o ? 7'b1000000 : 7'b1000001;
  /* fpu.vhdl:1745:17  */
  assign n16066_o = n16060_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:1732:17  */
  assign n16068_o = n16040_o ? n16048_o : 2'b00;
  /* fpu.vhdl:1732:17  */
  assign n16069_o = n16040_o ? n13151_o : n16063_o;
  /* fpu.vhdl:1732:17  */
  assign n16071_o = n16040_o & n16041_o;
  /* fpu.vhdl:1732:17  */
  assign n16073_o = n16040_o ? n16054_o : 1'b0;
  /* fpu.vhdl:1732:17  */
  assign n16075_o = n16040_o ? 1'b0 : n16066_o;
  /* fpu.vhdl:1732:17  */
  assign n16077_o = n16040_o ? n16057_o : 1'b0;
  /* fpu.vhdl:1730:13  */
  assign n16079_o = n13567_o == 7'b0100100;
  /* fpu.vhdl:1756:26  */
  assign n16081_o = r[21];
  /* fpu.vhdl:1756:30  */
  assign n16082_o = ~n16081_o;
  /* fpu.vhdl:1757:30  */
  assign n16083_o = r[20];
  /* fpu.vhdl:1757:34  */
  assign n16084_o = ~n16083_o;
  /* fpu.vhdl:1757:21  */
  assign n16087_o = n16084_o ? 7'b0100110 : 7'b0101110;
  /* fpu.vhdl:1762:29  */
  assign n16088_o = r[19];
  /* fpu.vhdl:1762:33  */
  assign n16089_o = ~n16088_o;
  /* fpu.vhdl:1762:17  */
  assign n16092_o = n16089_o ? 7'b0101011 : 7'b0101100;
  /* fpu.vhdl:1756:17  */
  assign n16093_o = n16082_o ? n16087_o : n16092_o;
  /* fpu.vhdl:1752:13  */
  assign n16095_o = n13567_o == 7'b0100101;
  /* fpu.vhdl:1773:22  */
  assign n16096_o = r[711:710];
  /* fpu.vhdl:1773:28  */
  assign n16098_o = n16096_o == 2'b00;
  /* fpu.vhdl:1773:17  */
  assign n16101_o = n16098_o ? 2'b01 : 2'b10;
  /* fpu.vhdl:1778:28  */
  assign n16102_o = r[709];
  /* fpu.vhdl:1780:42  */
  assign n16103_o = r[709];
  /* fpu.vhdl:1781:34  */
  assign n16104_o = multiply_to_f[0];
  /* fpu.vhdl:1783:34  */
  assign n16106_o = r[711:710];
  /* fpu.vhdl:1783:40  */
  assign n16108_o = n16106_o + 2'b01;
  assign n16110_o = {n16108_o, 1'b1};
  /* fpu.vhdl:1781:17  */
  assign n16111_o = n16104_o ? 7'b0100111 : n13151_o;
  assign n16112_o = {n13562_o, 1'b0};
  /* fpu.vhdl:1781:17  */
  assign n16113_o = n16104_o ? n16110_o : n16112_o;
  /* fpu.vhdl:1768:13  */
  assign n16115_o = n13567_o == 7'b0100110;
  /* fpu.vhdl:1791:42  */
  assign n16116_o = r[709];
  /* fpu.vhdl:1793:34  */
  assign n16117_o = multiply_to_f[0];
  /* fpu.vhdl:1795:26  */
  assign n16119_o = r[711:710];
  /* fpu.vhdl:1795:32  */
  assign n16121_o = n16119_o == 2'b11;
  /* fpu.vhdl:1795:21  */
  assign n16124_o = n16121_o ? 7'b0101000 : 7'b0100110;
  /* fpu.vhdl:1793:17  */
  assign n16125_o = n16117_o ? n16124_o : n13151_o;
  /* fpu.vhdl:1793:17  */
  assign n16126_o = n16117_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1787:13  */
  assign n16128_o = n13567_o == 7'b0100111;
  /* fpu.vhdl:1806:28  */
  assign n16129_o = r[709];
  /* fpu.vhdl:1807:42  */
  assign n16130_o = r[709];
  /* fpu.vhdl:1809:34  */
  assign n16131_o = multiply_to_f[0];
  /* fpu.vhdl:1809:17  */
  assign n16136_o = n16131_o ? 2'b10 : 2'b00;
  /* fpu.vhdl:1809:17  */
  assign n16137_o = n16131_o ? 7'b0101001 : n13151_o;
  /* fpu.vhdl:1809:17  */
  assign n16138_o = n16131_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1802:13  */
  assign n16140_o = n13567_o == 7'b0101000;
  /* fpu.vhdl:1821:42  */
  assign n16141_o = r[709];
  /* fpu.vhdl:1822:34  */
  assign n16142_o = multiply_to_f[0];
  /* fpu.vhdl:1822:17  */
  assign n16144_o = n16142_o ? 7'b0101010 : n13151_o;
  /* fpu.vhdl:1815:13  */
  assign n16146_o = n13567_o == 7'b0101001;
  /* fpu.vhdl:1830:31  */
  assign n16147_o = r[578];
  /* fpu.vhdl:1830:36  */
  assign n16148_o = n16147_o | n13538_o;
  /* fpu.vhdl:1834:28  */
  assign n16149_o = ~n13544_o;
  /* fpu.vhdl:1828:17  */
  assign n16152_o = n13551_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:1828:17  */
  assign n16153_o = n13551_o ? n16148_o : n16149_o;
  /* fpu.vhdl:1826:13  */
  assign n16156_o = n13567_o == 7'b0101010;
  /* fpu.vhdl:1838:13  */
  assign n16160_o = n13567_o == 7'b0101011;
  /* fpu.vhdl:1845:44  */
  assign n16161_o = n13530_o | n13535_o;
  /* fpu.vhdl:1846:35  */
  assign n16162_o = n13530_o | n13535_o;
  /* fpu.vhdl:1846:58  */
  assign n16163_o = r[238:159];
  /* fpu.vhdl:1846:60  */
  assign n16164_o = n16163_o[1:0];
  /* fpu.vhdl:1846:66  */
  assign n16166_o = n16164_o == 2'b00;
  /* fpu.vhdl:1846:53  */
  assign n16167_o = n16162_o | n16166_o;
  /* fpu.vhdl:1846:78  */
  assign n16168_o = r[709];
  /* fpu.vhdl:1846:84  */
  assign n16169_o = ~n16168_o;
  /* fpu.vhdl:1846:73  */
  assign n16170_o = n16167_o | n16169_o;
  /* fpu.vhdl:1850:34  */
  assign n16173_o = r[238:159];
  /* fpu.vhdl:1850:36  */
  assign n16174_o = n16173_o[15:3];
  /* fpu.vhdl:1846:17  */
  assign n16176_o = n16170_o ? 7'b0000000 : n13151_o;
  /* fpu.vhdl:1846:17  */
  assign n16177_o = n16170_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1846:17  */
  assign n16178_o = n16170_o ? 13'b0000000000000 : n16174_o;
  /* fpu.vhdl:1846:17  */
  assign n16179_o = n16170_o ? n13477_o : 2'b10;
  /* fpu.vhdl:1844:13  */
  assign n16181_o = n13567_o == 7'b0101101;
  /* fpu.vhdl:1857:41  */
  assign n16182_o = r[254];
  /* fpu.vhdl:1857:68  */
  assign n16183_o = r[254:243];
  /* fpu.vhdl:1857:54  */
  assign n16184_o = {n16182_o, n16183_o};
  /* fpu.vhdl:1858:33  */
  assign n16185_o = -n16184_o;
  /* fpu.vhdl:1854:13  */
  assign n16189_o = n13567_o == 7'b0101100;
  /* fpu.vhdl:1862:13  */
  assign n16195_o = n13567_o == 7'b0101110;
  /* fpu.vhdl:1875:13  */
  assign n16199_o = n13567_o == 7'b0101111;
  /* fpu.vhdl:1886:28  */
  assign n16200_o = r[709];
  /* fpu.vhdl:1888:34  */
  assign n16201_o = multiply_to_f[0];
  /* fpu.vhdl:1888:17  */
  assign n16206_o = n16201_o ? 2'b10 : 2'b00;
  /* fpu.vhdl:1888:17  */
  assign n16207_o = n16201_o ? 7'b0110001 : n13151_o;
  /* fpu.vhdl:1888:17  */
  assign n16208_o = n16201_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1883:13  */
  assign n16210_o = n13567_o == 7'b0110000;
  /* fpu.vhdl:1901:42  */
  assign n16211_o = r[709];
  /* fpu.vhdl:1903:34  */
  assign n16212_o = multiply_to_f[0];
  /* fpu.vhdl:1903:17  */
  assign n16214_o = n16212_o ? 7'b0110010 : n13151_o;
  /* fpu.vhdl:1895:13  */
  assign n16216_o = n13567_o == 7'b0110001;
  /* fpu.vhdl:1907:13  */
  assign n16221_o = n13567_o == 7'b0110010;
  /* fpu.vhdl:1919:42  */
  assign n16222_o = r[709];
  /* fpu.vhdl:1921:34  */
  assign n16223_o = multiply_to_f[0];
  /* fpu.vhdl:1921:17  */
  assign n16226_o = n16223_o ? 7'b0110100 : n13151_o;
  /* fpu.vhdl:1921:17  */
  assign n16227_o = n16223_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1915:13  */
  assign n16229_o = n13567_o == 7'b0110011;
  /* fpu.vhdl:1929:28  */
  assign n16230_o = r[709];
  /* fpu.vhdl:1932:34  */
  assign n16231_o = multiply_to_f[0];
  /* fpu.vhdl:1936:34  */
  assign n16233_o = r[711:710];
  /* fpu.vhdl:1936:40  */
  assign n16235_o = n16233_o + 2'b01;
  /* fpu.vhdl:1937:26  */
  assign n16236_o = r[711:710];
  /* fpu.vhdl:1937:32  */
  assign n16238_o = $unsigned(n16236_o) < $unsigned(2'b10);
  /* fpu.vhdl:1937:21  */
  assign n16242_o = n16238_o ? 7'b0110001 : 7'b0110101;
  /* fpu.vhdl:1937:21  */
  assign n16243_o = n16238_o ? 1'b1 : 1'b1;
  /* fpu.vhdl:1932:17  */
  assign n16246_o = n16231_o ? 2'b10 : 2'b00;
  assign n16247_o = {n16235_o, n16243_o};
  /* fpu.vhdl:1932:17  */
  assign n16248_o = n16231_o ? n16242_o : n13151_o;
  assign n16249_o = {n13562_o, 1'b0};
  /* fpu.vhdl:1932:17  */
  assign n16250_o = n16231_o ? n16247_o : n16249_o;
  /* fpu.vhdl:1926:13  */
  assign n16252_o = n13567_o == 7'b0110100;
  /* fpu.vhdl:1953:42  */
  assign n16253_o = r[709];
  /* fpu.vhdl:1954:34  */
  assign n16254_o = multiply_to_f[0];
  /* fpu.vhdl:1954:17  */
  assign n16257_o = n16254_o ? 7'b0110110 : n13151_o;
  /* fpu.vhdl:1954:17  */
  assign n16258_o = n16254_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:1945:13  */
  assign n16260_o = n13567_o == 7'b0110101;
  /* fpu.vhdl:1970:42  */
  assign n16261_o = r[709];
  /* fpu.vhdl:1971:34  */
  assign n16262_o = multiply_to_f[0];
  /* fpu.vhdl:1971:17  */
  assign n16264_o = n16262_o ? 7'b0110111 : n13151_o;
  /* fpu.vhdl:1959:13  */
  assign n16266_o = n13567_o == 7'b0110110;
  /* fpu.vhdl:1981:41  */
  assign n16267_o = r[254];
  /* fpu.vhdl:1981:68  */
  assign n16268_o = r[254:243];
  /* fpu.vhdl:1981:54  */
  assign n16269_o = {n16267_o, n16268_o};
  /* fpu.vhdl:1975:13  */
  assign n16274_o = n13567_o == 7'b0110111;
  /* fpu.vhdl:1994:42  */
  assign n16275_o = r[709];
  /* fpu.vhdl:1996:28  */
  assign n16276_o = r[709];
  /* fpu.vhdl:1997:34  */
  assign n16277_o = multiply_to_f[0];
  /* fpu.vhdl:1997:17  */
  assign n16279_o = n16277_o ? 7'b0111001 : n13151_o;
  /* fpu.vhdl:1987:13  */
  assign n16281_o = n13567_o == 7'b0111000;
  /* fpu.vhdl:2005:31  */
  assign n16282_o = r[578];
  /* fpu.vhdl:2005:36  */
  assign n16283_o = n16282_o | n13538_o;
  /* fpu.vhdl:2009:28  */
  assign n16284_o = ~n13544_o;
  /* fpu.vhdl:2003:17  */
  assign n16287_o = n13551_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:2003:17  */
  assign n16288_o = n13551_o ? n16283_o : n16284_o;
  /* fpu.vhdl:2001:13  */
  assign n16291_o = n13567_o == 7'b0111001;
  /* fpu.vhdl:2013:13  */
  assign n16295_o = n13567_o == 7'b0111010;
  /* fpu.vhdl:2023:40  */
  assign n16297_o = r[462:399];
  /* fpu.vhdl:2023:45  */
  assign n16298_o = r[519];
  /* fpu.vhdl:2023:55  */
  assign n16299_o = r[702:700];
  /* fpu.vhdl:2023:69  */
  assign n16300_o = r[648];
  /* fpu.vhdl:493:28  */
  assign n16308_o = n16297_o[1:0];
  /* fpu.vhdl:493:41  */
  assign n16309_o = {n16308_o, n16298_o};
  /* fpu.vhdl:494:28  */
  assign n16311_o = n16297_o[2];
  /* fpu.vhdl:500:19  */
  assign n16316_o = |(n16309_o);
  /* fpu.vhdl:501:16  */
  assign n16317_o = n16299_o[1:0];
  /* fpu.vhdl:503:24  */
  assign n16319_o = n16309_o == 3'b100;
  /* fpu.vhdl:503:38  */
  assign n16320_o = n16299_o[2];
  /* fpu.vhdl:503:42  */
  assign n16321_o = ~n16320_o;
  /* fpu.vhdl:503:32  */
  assign n16322_o = n16319_o & n16321_o;
  /* fpu.vhdl:506:34  */
  assign n16323_o = n16309_o[2];
  /* fpu.vhdl:503:17  */
  assign n16324_o = n16322_o ? n16311_o : n16323_o;
  /* fpu.vhdl:502:13  */
  assign n16326_o = n16317_o == 2'b00;
  /* fpu.vhdl:508:13  */
  assign n16328_o = n16317_o == 2'b01;
  /* fpu.vhdl:510:22  */
  assign n16329_o = n16299_o[0];
  /* fpu.vhdl:510:26  */
  assign n16330_o = n16329_o == n16300_o;
  assign n16331_o = {1'b0, n16316_o};
  /* fpu.vhdl:512:34  */
  assign n16332_o = n16331_o[0];
  /* fpu.vhdl:510:17  */
  assign n16333_o = n16330_o ? n16332_o : 1'b0;
  assign n16334_o = {n16328_o, n16326_o};
  /* fpu.vhdl:501:9  */
  always @*
    case (n16334_o)
      2'b10: n16335_o = 1'b0;
      2'b01: n16335_o = n16324_o;
      default: n16335_o = n16333_o;
    endcase
  assign n16336_o = {n16335_o, n16316_o};
  /* fpu.vhdl:2026:26  */
  assign n16337_o = r[25];
  /* fpu.vhdl:2026:42  */
  assign n16338_o = r[648];
  /* fpu.vhdl:2026:36  */
  assign n16339_o = n16337_o & n16338_o;
  /* fpu.vhdl:2027:30  */
  assign n16340_o = r_hi_nz | r_lo_nz;
  assign n16341_o = r[143:127];
  assign n16342_o = r[158:146];
  assign n16343_o = {n13479_o, n13564_o, 2'b00, n13477_o, n13562_o, 1'b0, n13475_o, 1'b0, n13558_o, n13473_o, n13487_o, n13471_o, 1'b0, 13'b0000000000000, n13560_o, n13469_o, n16342_o, n16336_o, n16341_o, n13467_o, n13556_o, 1'b0, 1'b0, n13151_o};
  /* fpu.vhdl:2027:51  */
  assign n16344_o = n16343_o[145];
  /* fpu.vhdl:2027:41  */
  assign n16345_o = n16340_o | n16344_o;
  /* fpu.vhdl:2026:60  */
  assign n16346_o = n16339_o & n16345_o;
  /* fpu.vhdl:2026:17  */
  assign n16349_o = n16346_o ? 7'b0111111 : 7'b0111101;
  /* fpu.vhdl:2020:13  */
  assign n16351_o = n13567_o == 7'b0111011;
  /* fpu.vhdl:2033:13  */
  assign n16354_o = n13567_o == 7'b0111100;
  /* fpu.vhdl:2040:33  */
  assign n16355_o = r[648];
  /* fpu.vhdl:2041:36  */
  assign n16356_o = r[145];
  /* fpu.vhdl:2041:53  */
  assign n16357_o = r[648];
  /* fpu.vhdl:2041:47  */
  assign n16358_o = n16356_o ^ n16357_o;
  /* fpu.vhdl:2043:28  */
  assign n16359_o = r[26:25];
  /* fpu.vhdl:2045:42  */
  assign n16360_o = r[430];
  /* fpu.vhdl:2045:54  */
  assign n16361_o = r[429];
  /* fpu.vhdl:2045:69  */
  assign n16362_o = r[648];
  /* fpu.vhdl:2045:63  */
  assign n16363_o = ~n16362_o;
  /* fpu.vhdl:2045:59  */
  assign n16364_o = n16361_o & n16363_o;
  /* fpu.vhdl:2045:47  */
  assign n16365_o = n16360_o | n16364_o;
  /* fpu.vhdl:2044:21  */
  assign n16367_o = n16359_o == 2'b00;
  /* fpu.vhdl:2047:42  */
  assign n16368_o = r[430];
  /* fpu.vhdl:2046:21  */
  assign n16370_o = n16359_o == 2'b01;
  /* fpu.vhdl:2049:42  */
  assign n16371_o = r[462];
  /* fpu.vhdl:2049:54  */
  assign n16372_o = r[461];
  /* fpu.vhdl:2049:69  */
  assign n16373_o = r[648];
  /* fpu.vhdl:2049:63  */
  assign n16374_o = ~n16373_o;
  /* fpu.vhdl:2049:59  */
  assign n16375_o = n16372_o & n16374_o;
  /* fpu.vhdl:2049:47  */
  assign n16376_o = n16371_o | n16375_o;
  /* fpu.vhdl:2048:21  */
  assign n16378_o = n16359_o == 2'b10;
  /* fpu.vhdl:2051:42  */
  assign n16379_o = r[462];
  assign n16380_o = {n16378_o, n16370_o, n16367_o};
  /* fpu.vhdl:2043:17  */
  always @*
    case (n16380_o)
      3'b100: n16381_o = n16376_o;
      3'b010: n16381_o = n16368_o;
      3'b001: n16381_o = n16365_o;
      default: n16381_o = n16379_o;
    endcase
  /* fpu.vhdl:2056:31  */
  assign n16383_o = r[144];
  assign n16385_o = r[152];
  /* fpu.vhdl:2056:21  */
  assign n16386_o = n16383_o ? 1'b1 : n16385_o;
  /* fpu.vhdl:2053:17  */
  assign n16387_o = n16381_o ? 7'b0111110 : n13151_o;
  assign n16388_o = r[152];
  /* fpu.vhdl:2053:17  */
  assign n16389_o = n16381_o ? n16388_o : n16386_o;
  /* fpu.vhdl:2053:17  */
  assign n16392_o = n16381_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:2038:13  */
  assign n16394_o = n13567_o == 7'b0111101;
  /* fpu.vhdl:2063:26  */
  assign n16395_o = r[26];
  /* fpu.vhdl:2063:30  */
  assign n16396_o = ~n16395_o;
  /* fpu.vhdl:2064:31  */
  assign n16397_o = r[430];
  /* fpu.vhdl:2066:31  */
  assign n16398_o = r[462];
  /* fpu.vhdl:2063:17  */
  assign n16399_o = n16396_o ? n16397_o : n16398_o;
  /* fpu.vhdl:2068:41  */
  assign n16400_o = r[26:25];
  /* fpu.vhdl:2068:33  */
  assign n16402_o = {1'b1, n16400_o};
  /* fpu.vhdl:2068:58  */
  assign n16403_o = r[648];
  /* fpu.vhdl:2068:54  */
  assign n16404_o = {n16402_o, n16403_o};
  /* fpu.vhdl:2069:27  */
  assign n16405_o = r[25];
  /* fpu.vhdl:2069:31  */
  assign n16406_o = ~n16405_o;
  /* fpu.vhdl:2069:50  */
  assign n16407_o = r[648];
  /* fpu.vhdl:2069:45  */
  assign n16408_o = n16399_o != n16407_o;
  /* fpu.vhdl:2069:37  */
  assign n16409_o = n16406_o & n16408_o;
  /* fpu.vhdl:2070:28  */
  assign n16410_o = r[25];
  /* fpu.vhdl:2070:46  */
  assign n16412_o = n16399_o != 1'b1;
  /* fpu.vhdl:2070:38  */
  assign n16413_o = n16410_o & n16412_o;
  /* fpu.vhdl:2069:63  */
  assign n16414_o = n16409_o | n16413_o;
  /* fpu.vhdl:2075:31  */
  assign n16416_o = r[144];
  assign n16418_o = r[152];
  /* fpu.vhdl:2075:21  */
  assign n16419_o = n16416_o ? 1'b1 : n16418_o;
  /* fpu.vhdl:2069:17  */
  assign n16422_o = n16414_o ? 2'b11 : 2'b00;
  assign n16423_o = r[135];
  /* fpu.vhdl:2069:17  */
  assign n16424_o = n16414_o ? 1'b1 : n16423_o;
  assign n16425_o = r[152];
  /* fpu.vhdl:2069:17  */
  assign n16426_o = n16414_o ? n16425_o : n16419_o;
  /* fpu.vhdl:2069:17  */
  assign n16429_o = n16414_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:2062:13  */
  assign n16431_o = n13567_o == 7'b0111110;
  /* fpu.vhdl:2083:41  */
  assign n16432_o = r[26:25];
  /* fpu.vhdl:2083:33  */
  assign n16434_o = {1'b1, n16432_o};
  /* fpu.vhdl:2083:58  */
  assign n16435_o = r[648];
  /* fpu.vhdl:2083:54  */
  assign n16436_o = {n16434_o, n16435_o};
  /* fpu.vhdl:2084:22  */
  assign n16437_o = r[318:239];
  /* fpu.vhdl:2084:24  */
  assign n16438_o = n16437_o[1:0];
  /* fpu.vhdl:2084:30  */
  assign n16440_o = n16438_o == 2'b11;
  assign n16442_o = n16436_o[0];
  /* fpu.vhdl:2084:17  */
  assign n16443_o = n16440_o ? 1'b1 : n16442_o;
  assign n16444_o = n16436_o[3:1];
  /* fpu.vhdl:2081:13  */
  assign n16447_o = n13567_o == 7'b0111111;
  /* fpu.vhdl:2091:13  */
  assign n16450_o = n13567_o == 7'b0010111;
  /* fpu.vhdl:2098:22  */
  assign n16451_o = r[707];
  /* fpu.vhdl:2098:40  */
  assign n16452_o = n16451_o & n13538_o;
  assign n16454_o = r[519];
  /* fpu.vhdl:2098:17  */
  assign n16455_o = n16452_o ? 1'b1 : n16454_o;
  /* fpu.vhdl:2101:23  */
  assign n16456_o = r[462:453];
  /* fpu.vhdl:2101:38  */
  assign n16458_o = n16456_o != 10'b0000000001;
  /* fpu.vhdl:2107:44  */
  assign n16460_o = n13526_o - n13518_o;
  /* fpu.vhdl:2109:21  */
  assign n16464_o = n13535_o ? 7'b1000011 : 7'b1000100;
  /* fpu.vhdl:2106:21  */
  assign n16465_o = n13530_o ? 7'b1000010 : n16464_o;
  /* fpu.vhdl:2106:21  */
  assign n16466_o = n13530_o ? n16460_o : 13'b0000000000000;
  /* fpu.vhdl:2101:17  */
  assign n16467_o = n16458_o ? 7'b1000001 : n16465_o;
  /* fpu.vhdl:2101:17  */
  assign n16468_o = n16458_o ? 13'b0000000000000 : n16466_o;
  /* fpu.vhdl:2101:17  */
  assign n16471_o = n16458_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:2101:17  */
  assign n16474_o = n16458_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:2097:13  */
  assign n16476_o = n13567_o == 7'b1000000;
  /* fpu.vhdl:2122:40  */
  assign n16477_o = n13526_o - n13518_o;
  /* fpu.vhdl:2124:17  */
  assign n16481_o = n13535_o ? 7'b1000011 : 7'b1000100;
  /* fpu.vhdl:2121:17  */
  assign n16482_o = n13530_o ? 7'b1000010 : n16481_o;
  /* fpu.vhdl:2121:17  */
  assign n16483_o = n13530_o ? n16477_o : 13'b0000000000000;
  /* fpu.vhdl:2116:13  */
  assign n16485_o = n13567_o == 7'b1000001;
  /* fpu.vhdl:2133:27  */
  assign n16487_o = r[132];
  /* fpu.vhdl:2133:38  */
  assign n16488_o = ~n16487_o;
  /* fpu.vhdl:2143:39  */
  assign n16491_o = r[663:651];
  /* fpu.vhdl:2143:50  */
  assign n16492_o = n16491_o + n13523_o;
  /* fpu.vhdl:2144:27  */
  assign n16493_o = r[453];
  /* fpu.vhdl:2144:32  */
  assign n16494_o = ~n16493_o;
  /* fpu.vhdl:2144:21  */
  assign n16497_o = n16494_o ? 7'b1000001 : 7'b1000100;
  /* fpu.vhdl:2144:21  */
  assign n16500_o = n16494_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:2133:17  */
  assign n16503_o = n16488_o ? 2'b01 : 2'b00;
  /* fpu.vhdl:2133:17  */
  assign n16504_o = n16488_o ? 7'b1000100 : n16497_o;
  assign n16505_o = r[154];
  /* fpu.vhdl:2133:17  */
  assign n16506_o = n16488_o ? n16505_o : 1'b1;
  assign n16507_o = r[663:651];
  /* fpu.vhdl:2133:17  */
  assign n16508_o = n16488_o ? n16507_o : n16492_o;
  /* fpu.vhdl:2133:17  */
  assign n16510_o = n16488_o ? 1'b0 : n16500_o;
  /* fpu.vhdl:2133:17  */
  assign n16513_o = n16488_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:2130:13  */
  assign n16515_o = n13567_o == 7'b1000010;
  /* fpu.vhdl:2154:27  */
  assign n16517_o = r[133];
  /* fpu.vhdl:2154:38  */
  assign n16518_o = ~n16517_o;
  /* fpu.vhdl:2159:36  */
  assign n16521_o = r[701:700];
  /* fpu.vhdl:2159:49  */
  assign n16523_o = n16521_o == 2'b00;
  /* fpu.vhdl:2160:38  */
  assign n16524_o = r[701];
  /* fpu.vhdl:2160:64  */
  assign n16525_o = r[700];
  /* fpu.vhdl:2160:72  */
  assign n16526_o = r[648];
  /* fpu.vhdl:2160:68  */
  assign n16527_o = n16525_o == n16526_o;
  /* fpu.vhdl:2160:48  */
  assign n16528_o = n16524_o & n16527_o;
  /* fpu.vhdl:2159:56  */
  assign n16529_o = n16523_o | n16528_o;
  /* fpu.vhdl:2159:21  */
  assign n16533_o = n16529_o ? 1'b1 : 1'b0;
  assign n16534_o = r[650:649];
  /* fpu.vhdl:2159:21  */
  assign n16535_o = n16529_o ? 2'b10 : n16534_o;
  /* fpu.vhdl:2169:43  */
  assign n16536_o = r[126];
  /* fpu.vhdl:2169:39  */
  assign n16538_o = {3'b001, n16536_o};
  /* fpu.vhdl:2173:39  */
  assign n16539_o = r[663:651];
  /* fpu.vhdl:2173:50  */
  assign n16540_o = n16539_o - n13523_o;
  /* fpu.vhdl:2154:17  */
  assign n16544_o = n16518_o ? 2'b11 : 2'b00;
  /* fpu.vhdl:2154:17  */
  assign n16546_o = n16518_o ? n16538_o : 4'b0000;
  assign n16547_o = {n16533_o, 1'b1};
  assign n16548_o = {n13520_o, n16535_o};
  /* fpu.vhdl:2154:17  */
  assign n16549_o = n16518_o ? n13151_o : 7'b1000100;
  assign n16550_o = r[145:144];
  /* fpu.vhdl:2154:17  */
  assign n16551_o = n16518_o ? n16547_o : n16550_o;
  assign n16552_o = r[152];
  /* fpu.vhdl:2154:17  */
  assign n16553_o = n16518_o ? 1'b1 : n16552_o;
  assign n16554_o = n16548_o[1:0];
  assign n16555_o = r[650:649];
  /* fpu.vhdl:2154:17  */
  assign n16556_o = n16518_o ? n16554_o : n16555_o;
  assign n16557_o = n16548_o[14:2];
  /* fpu.vhdl:2154:17  */
  assign n16558_o = n16518_o ? n16557_o : n16540_o;
  /* fpu.vhdl:2154:17  */
  assign n16561_o = n16518_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:2152:13  */
  assign n16563_o = n13567_o == 7'b1000011;
  /* fpu.vhdl:2179:40  */
  assign n16565_o = r[462:399];
  /* fpu.vhdl:2179:45  */
  assign n16566_o = r[519];
  /* fpu.vhdl:2179:50  */
  assign n16567_o = r[126];
  /* fpu.vhdl:2179:65  */
  assign n16568_o = r[702:700];
  /* fpu.vhdl:2179:79  */
  assign n16569_o = r[648];
  /* fpu.vhdl:492:24  */
  assign n16577_o = ~n16567_o;
  /* fpu.vhdl:493:28  */
  assign n16578_o = n16565_o[1:0];
  /* fpu.vhdl:493:41  */
  assign n16579_o = {n16578_o, n16566_o};
  /* fpu.vhdl:494:28  */
  assign n16580_o = n16565_o[2];
  /* fpu.vhdl:496:28  */
  assign n16581_o = n16565_o[30:29];
  /* fpu.vhdl:496:43  */
  assign n16582_o = {n16581_o, n16566_o};
  /* fpu.vhdl:497:28  */
  assign n16583_o = n16565_o[31];
  /* fpu.vhdl:492:9  */
  assign n16584_o = n16577_o ? n16579_o : n16582_o;
  /* fpu.vhdl:492:9  */
  assign n16586_o = n16577_o ? n16580_o : n16583_o;
  /* fpu.vhdl:500:19  */
  assign n16591_o = |(n16584_o);
  /* fpu.vhdl:501:16  */
  assign n16592_o = n16568_o[1:0];
  /* fpu.vhdl:503:24  */
  assign n16594_o = n16584_o == 3'b100;
  /* fpu.vhdl:503:38  */
  assign n16595_o = n16568_o[2];
  /* fpu.vhdl:503:42  */
  assign n16596_o = ~n16595_o;
  /* fpu.vhdl:503:32  */
  assign n16597_o = n16594_o & n16596_o;
  /* fpu.vhdl:506:34  */
  assign n16598_o = n16584_o[2];
  /* fpu.vhdl:503:17  */
  assign n16599_o = n16597_o ? n16586_o : n16598_o;
  /* fpu.vhdl:502:13  */
  assign n16601_o = n16592_o == 2'b00;
  /* fpu.vhdl:508:13  */
  assign n16603_o = n16592_o == 2'b01;
  /* fpu.vhdl:510:22  */
  assign n16604_o = n16568_o[0];
  /* fpu.vhdl:510:26  */
  assign n16605_o = n16604_o == n16569_o;
  assign n16606_o = {1'b0, n16591_o};
  /* fpu.vhdl:512:34  */
  assign n16607_o = n16606_o[0];
  /* fpu.vhdl:510:17  */
  assign n16608_o = n16605_o ? n16607_o : 1'b0;
  assign n16609_o = {n16603_o, n16601_o};
  /* fpu.vhdl:501:9  */
  always @*
    case (n16609_o)
      2'b10: n16610_o = 1'b0;
      2'b01: n16610_o = n16599_o;
      default: n16610_o = n16608_o;
    endcase
  assign n16611_o = {n16610_o, n16591_o};
  /* fpu.vhdl:2181:25  */
  assign n16612_o = n16611_o[1];
  /* fpu.vhdl:2187:27  */
  assign n16615_o = r[453];
  /* fpu.vhdl:2187:32  */
  assign n16616_o = ~n16615_o;
  /* fpu.vhdl:2187:21  */
  assign n16618_o = n16616_o ? 7'b1000110 : n13151_o;
  /* fpu.vhdl:2187:21  */
  assign n16621_o = n16616_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:2187:21  */
  assign n16624_o = n16616_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:2181:17  */
  assign n16627_o = n16612_o ? 2'b10 : 2'b00;
  /* fpu.vhdl:2181:17  */
  assign n16628_o = n16612_o ? 7'b1000101 : n16618_o;
  /* fpu.vhdl:2181:17  */
  assign n16629_o = n16612_o ? 13'b1111111111111 : 13'b0000000000000;
  /* fpu.vhdl:2181:17  */
  assign n16631_o = n16612_o ? 1'b0 : n16621_o;
  /* fpu.vhdl:2181:17  */
  assign n16633_o = n16612_o ? 1'b0 : n16624_o;
  /* fpu.vhdl:2196:25  */
  assign n16634_o = n16611_o[0];
  /* fpu.vhdl:2198:26  */
  assign n16636_o = r[698];
  assign n16638_o = r[154];
  /* fpu.vhdl:2196:17  */
  assign n16639_o = n16643_o ? 1'b1 : n16638_o;
  assign n16640_o = r[152];
  /* fpu.vhdl:2196:17  */
  assign n16641_o = n16634_o ? 1'b1 : n16640_o;
  /* fpu.vhdl:2196:17  */
  assign n16643_o = n16634_o & n16636_o;
  /* fpu.vhdl:2177:13  */
  assign n16645_o = n13567_o == 7'b1000100;
  /* fpu.vhdl:2207:23  */
  assign n16647_o = r[454];
  /* fpu.vhdl:2209:21  */
  assign n16649_o = n13535_o ? 7'b1000011 : n13151_o;
  /* fpu.vhdl:2209:21  */
  assign n16652_o = n13535_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:2214:26  */
  assign n16653_o = r[453];
  /* fpu.vhdl:2214:31  */
  assign n16654_o = ~n16653_o;
  /* fpu.vhdl:2214:17  */
  assign n16656_o = n16654_o ? 7'b1000110 : n13151_o;
  /* fpu.vhdl:2214:17  */
  assign n16659_o = n16654_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:2214:17  */
  assign n16662_o = n16654_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:2207:17  */
  assign n16665_o = n16647_o ? 2'b01 : 2'b00;
  /* fpu.vhdl:2207:17  */
  assign n16666_o = n16647_o ? n16649_o : n16656_o;
  /* fpu.vhdl:2207:17  */
  assign n16667_o = n16647_o ? n16652_o : n16659_o;
  /* fpu.vhdl:2207:17  */
  assign n16669_o = n16647_o ? 1'b0 : n16662_o;
  /* fpu.vhdl:2203:13  */
  assign n16671_o = n13567_o == 7'b1000101;
  /* fpu.vhdl:2224:58  */
  assign n16672_o = r[126];
  /* fpu.vhdl:2224:52  */
  assign n16673_o = ~n16672_o;
  /* fpu.vhdl:2224:48  */
  assign n16674_o = r_lo_nz & n16673_o;
  /* fpu.vhdl:2224:36  */
  assign n16675_o = r_hi_nz | n16674_o;
  /* fpu.vhdl:2225:28  */
  assign n16676_o = ~n16675_o;
  /* fpu.vhdl:2227:26  */
  assign n16678_o = r[703];
  /* fpu.vhdl:2229:54  */
  assign n16679_o = r[701];
  /* fpu.vhdl:2229:74  */
  assign n16680_o = r[700];
  /* fpu.vhdl:2229:58  */
  assign n16681_o = n16679_o & n16680_o;
  assign n16682_o = r[648];
  /* fpu.vhdl:2227:21  */
  assign n16683_o = n16678_o ? n16681_o : n16682_o;
  /* fpu.vhdl:2236:40  */
  assign n16685_o = n13526_o - 13'b1110000000010;
  /* fpu.vhdl:2237:32  */
  assign n16687_o = $signed(n13526_o) < $signed(13'b1110000000010);
  /* fpu.vhdl:2237:21  */
  assign n16689_o = n16687_o ? 7'b1000111 : n13151_o;
  /* fpu.vhdl:2237:21  */
  assign n16692_o = n16687_o ? 1'b0 : 1'b1;
  /* fpu.vhdl:2225:17  */
  assign n16695_o = n16676_o ? 2'b00 : 2'b01;
  assign n16696_o = {2'b00, n16683_o};
  /* fpu.vhdl:2225:17  */
  assign n16697_o = n16676_o ? n13151_o : n16689_o;
  assign n16698_o = r[650:648];
  /* fpu.vhdl:2225:17  */
  assign n16699_o = n16676_o ? n16696_o : n16698_o;
  /* fpu.vhdl:2225:17  */
  assign n16700_o = n16676_o ? 13'b0000000000000 : n16685_o;
  assign n16701_o = n13465_o[2];
  assign n16702_o = r[699];
  /* fpu.vhdl:650:9  */
  assign n16703_o = n13152_o ? n16701_o : n16702_o;
  /* fpu.vhdl:2225:17  */
  assign n16704_o = n16676_o ? n16703_o : n13530_o;
  /* fpu.vhdl:2225:17  */
  assign n16706_o = n16676_o ? 1'b1 : n16692_o;
  /* fpu.vhdl:2222:13  */
  assign n16708_o = n13567_o == 7'b1000110;
  /* fpu.vhdl:2244:13  */
  assign n16710_o = n13567_o == 7'b1000111;
  /* fpu.vhdl:2250:23  */
  assign n16711_o = r[716];
  /* fpu.vhdl:2250:41  */
  assign n16712_o = r[238:159];
  /* fpu.vhdl:2250:43  */
  assign n16713_o = n16712_o[1:0];
  /* fpu.vhdl:2250:49  */
  assign n16715_o = n16713_o == 2'b11;
  /* fpu.vhdl:2250:35  */
  assign n16716_o = n16711_o & n16715_o;
  /* fpu.vhdl:2250:71  */
  assign n16717_o = r[228];
  /* fpu.vhdl:2250:76  */
  assign n16718_o = ~n16717_o;
  /* fpu.vhdl:2250:55  */
  assign n16719_o = n16716_o & n16718_o;
  /* fpu.vhdl:2251:24  */
  assign n16720_o = r[717];
  /* fpu.vhdl:2251:42  */
  assign n16721_o = r[318:239];
  /* fpu.vhdl:2251:44  */
  assign n16722_o = n16721_o[1:0];
  /* fpu.vhdl:2251:50  */
  assign n16724_o = n16722_o == 2'b11;
  /* fpu.vhdl:2251:36  */
  assign n16725_o = n16720_o & n16724_o;
  /* fpu.vhdl:2251:72  */
  assign n16726_o = r[308];
  /* fpu.vhdl:2251:77  */
  assign n16727_o = ~n16726_o;
  /* fpu.vhdl:2251:56  */
  assign n16728_o = n16725_o & n16727_o;
  /* fpu.vhdl:2250:83  */
  assign n16729_o = n16719_o | n16728_o;
  /* fpu.vhdl:2252:24  */
  assign n16730_o = r[718];
  /* fpu.vhdl:2252:42  */
  assign n16731_o = r[398:319];
  /* fpu.vhdl:2252:44  */
  assign n16732_o = n16731_o[1:0];
  /* fpu.vhdl:2252:50  */
  assign n16734_o = n16732_o == 2'b11;
  /* fpu.vhdl:2252:36  */
  assign n16735_o = n16730_o & n16734_o;
  /* fpu.vhdl:2252:72  */
  assign n16736_o = r[388];
  /* fpu.vhdl:2252:77  */
  assign n16737_o = ~n16736_o;
  /* fpu.vhdl:2252:56  */
  assign n16738_o = n16735_o & n16737_o;
  /* fpu.vhdl:2251:84  */
  assign n16739_o = n16729_o | n16738_o;
  assign n16741_o = r[151];
  /* fpu.vhdl:2250:17  */
  assign n16742_o = n16739_o ? 1'b1 : n16741_o;
  /* fpu.vhdl:2250:17  */
  assign n16745_o = n16739_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:2257:22  */
  assign n16746_o = r[716];
  /* fpu.vhdl:2257:40  */
  assign n16747_o = r[238:159];
  /* fpu.vhdl:2257:42  */
  assign n16748_o = n16747_o[1:0];
  /* fpu.vhdl:2257:48  */
  assign n16750_o = n16748_o == 2'b11;
  /* fpu.vhdl:2257:34  */
  assign n16751_o = n16746_o & n16750_o;
  /* fpu.vhdl:2259:25  */
  assign n16753_o = r[717];
  /* fpu.vhdl:2259:43  */
  assign n16754_o = r[318:239];
  /* fpu.vhdl:2259:45  */
  assign n16755_o = n16754_o[1:0];
  /* fpu.vhdl:2259:51  */
  assign n16757_o = n16755_o == 2'b11;
  /* fpu.vhdl:2259:37  */
  assign n16758_o = n16753_o & n16757_o;
  /* fpu.vhdl:2261:25  */
  assign n16760_o = r[718];
  /* fpu.vhdl:2261:43  */
  assign n16761_o = r[398:319];
  /* fpu.vhdl:2261:45  */
  assign n16762_o = n16761_o[1:0];
  /* fpu.vhdl:2261:51  */
  assign n16764_o = n16762_o == 2'b11;
  /* fpu.vhdl:2261:37  */
  assign n16765_o = n16760_o & n16764_o;
  /* fpu.vhdl:2261:17  */
  assign n16767_o = n16765_o ? 2'b11 : 2'b00;
  /* fpu.vhdl:2259:17  */
  assign n16768_o = n16758_o ? 2'b10 : n16767_o;
  /* fpu.vhdl:2257:17  */
  assign n16769_o = n16751_o ? 2'b01 : n16768_o;
  /* fpu.vhdl:2249:13  */
  assign n16772_o = n13567_o == 7'b1001110;
  /* fpu.vhdl:2268:24  */
  assign n16773_o = r[715:714];
  /* fpu.vhdl:2270:44  */
  assign n16774_o = r[318:239];
  /* fpu.vhdl:2270:46  */
  assign n16775_o = n16774_o[2];
  /* fpu.vhdl:2270:61  */
  assign n16776_o = r[720];
  /* fpu.vhdl:2270:55  */
  assign n16777_o = n16775_o ^ n16776_o;
  /* fpu.vhdl:2271:43  */
  assign n16778_o = r[318:239];
  /* fpu.vhdl:2271:45  */
  assign n16779_o = n16778_o[15:3];
  /* fpu.vhdl:2272:45  */
  assign n16780_o = r[318:239];
  /* fpu.vhdl:2272:47  */
  assign n16781_o = n16780_o[1:0];
  /* fpu.vhdl:2269:21  */
  assign n16783_o = n16773_o == 2'b10;
  /* fpu.vhdl:2274:44  */
  assign n16784_o = r[398:319];
  /* fpu.vhdl:2274:46  */
  assign n16785_o = n16784_o[2];
  /* fpu.vhdl:2274:61  */
  assign n16786_o = r[720];
  /* fpu.vhdl:2274:55  */
  assign n16787_o = n16785_o ^ n16786_o;
  /* fpu.vhdl:2275:43  */
  assign n16788_o = r[398:319];
  /* fpu.vhdl:2275:45  */
  assign n16789_o = n16788_o[15:3];
  /* fpu.vhdl:2276:45  */
  assign n16790_o = r[398:319];
  /* fpu.vhdl:2276:47  */
  assign n16791_o = n16790_o[1:0];
  /* fpu.vhdl:2273:21  */
  assign n16793_o = n16773_o == 2'b11;
  /* fpu.vhdl:2278:44  */
  assign n16794_o = r[238:159];
  /* fpu.vhdl:2278:46  */
  assign n16795_o = n16794_o[2];
  /* fpu.vhdl:2278:61  */
  assign n16796_o = r[720];
  /* fpu.vhdl:2278:55  */
  assign n16797_o = n16795_o ^ n16796_o;
  /* fpu.vhdl:2279:43  */
  assign n16798_o = r[238:159];
  /* fpu.vhdl:2279:45  */
  assign n16799_o = n16798_o[15:3];
  /* fpu.vhdl:2280:45  */
  assign n16800_o = r[238:159];
  /* fpu.vhdl:2280:47  */
  assign n16801_o = n16800_o[1:0];
  assign n16802_o = {n16793_o, n16783_o};
  /* fpu.vhdl:2268:17  */
  always @*
    case (n16802_o)
      2'b10: n16803_o = n16787_o;
      2'b01: n16803_o = n16777_o;
      default: n16803_o = n16797_o;
    endcase
  /* fpu.vhdl:2268:17  */
  always @*
    case (n16802_o)
      2'b10: n16804_o = n16791_o;
      2'b01: n16804_o = n16781_o;
      default: n16804_o = n16801_o;
    endcase
  /* fpu.vhdl:2268:17  */
  always @*
    case (n16802_o)
      2'b10: n16805_o = n16789_o;
      2'b01: n16805_o = n16779_o;
      default: n16805_o = n16799_o;
    endcase
  /* fpu.vhdl:2266:13  */
  assign n16807_o = n13567_o == 7'b1001111;
  assign n16808_o = {n16807_o, n16772_o, n16710_o, n16708_o, n16671_o, n16645_o, n16563_o, n16515_o, n16485_o, n16476_o, n16450_o, n16447_o, n16431_o, n16394_o, n16354_o, n16351_o, n16295_o, n16291_o, n16281_o, n16274_o, n16266_o, n16260_o, n16252_o, n16229_o, n16221_o, n16216_o, n16210_o, n16199_o, n16195_o, n16189_o, n16181_o, n16160_o, n16156_o, n16146_o, n16140_o, n16128_o, n16115_o, n16095_o, n16079_o, n16032_o, n16009_o, n16002_o, n15998_o, n15992_o, n15973_o, n15967_o, n15939_o, n15936_o, n15858_o, n15849_o, n15841_o, n15830_o, n15802_o, n15799_o, n15789_o, n15785_o, n15734_o, n15727_o, n15440_o, n15365_o, n15318_o, n15247_o, n15225_o, n15096_o, n14973_o, n14809_o, n14779_o, n14697_o, n14647_o, n14591_o, n14564_o, n14521_o, n14482_o, n14471_o, n14349_o, n14176_o, n13972_o, n13919_o, n13841_o, n13751_o};
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16814_o = n16627_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b11;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16814_o = 2'b01;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16814_o = 2'b01;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16814_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16814_o = 2'b00;
      default: n16814_o = 2'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b01;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16836_o = n16695_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16836_o = n16665_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16836_o = n16544_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16836_o = n16503_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b01;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b01;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b11;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16836_o = n16422_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b01;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b01;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b01;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16836_o = n16246_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16836_o = n16206_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16836_o = 2'b01;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16836_o = 2'b11;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16836_o = 2'b11;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16836_o = 2'b11;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16836_o = n16136_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16836_o = n16068_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16836_o = 2'b10;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16836_o = 2'b01;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16836_o = 2'b10;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16836_o = 2'b10;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16836_o = n15916_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16836_o = 2'b01;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16836_o = 2'b11;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16836_o = 2'b11;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16836_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16836_o = 2'b00;
      default: n16836_o = 2'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16843_o = n16018_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16843_o = 2'b11;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16843_o = 2'b10;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16843_o = 2'b11;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16843_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16843_o = 2'b00;
      default: n16843_o = 2'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16847_o = n16355_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16847_o = n16021_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16847_o = n15919_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16847_o = n14789_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16847_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16847_o = 1'b0;
      default: n16847_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b1;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16852_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16852_o = 1'b0;
      default: n16852_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16857_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16857_o = n15850_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16857_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16857_o = 1'b0;
      default: n16857_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16862_o = n16358_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16862_o = n16287_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16862_o = n16152_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16862_o = n16023_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16862_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16862_o = n15922_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16862_o = n15854_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16862_o = n14792_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16862_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16862_o = 1'b0;
      default: n16862_o = 1'bX;
    endcase
  assign n16864_o = n14476_o[0];
  assign n16868_o = n16404_o[0];
  assign n16869_o = n16546_o[0];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16872_o = n16869_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16872_o = n16443_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16872_o = n16868_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16872_o = 1'b1;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16872_o = 1'b1;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16872_o = 1'b1;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16872_o = n16864_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16872_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16872_o = 1'b0;
      default: n16872_o = 1'bX;
    endcase
  assign n16873_o = n14476_o[3:1];
  assign n16877_o = n16404_o[3:1];
  assign n16878_o = n16546_o[3:1];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16881_o = n16878_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16881_o = n16444_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16881_o = n16877_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16881_o = 3'b011;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16881_o = 3'b011;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16881_o = 3'b011;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16881_o = n16873_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16881_o = 3'b000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16881_o = 3'b000;
      default: n16881_o = 3'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16885_o = n16275_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16885_o = n16261_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16885_o = n16253_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16885_o = n16222_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16885_o = 1'b1;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16885_o = n16211_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16885_o = 1'b1;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16885_o = n16141_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16885_o = n16130_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16885_o = n16116_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16885_o = n16103_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16885_o = n16003_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16885_o = n15985_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16885_o = n15968_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16885_o = n15698_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16885_o = n15082_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16885_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16885_o = 1'b0;
      default: n16885_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b11;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b10;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b11;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16899_o = 2'b11;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16899_o = 2'b10;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16899_o = 2'b10;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16899_o = 2'b01;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16899_o = 2'b01;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16899_o = 2'b10;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16899_o = 2'b01;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16899_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16899_o = 2'b00;
      default: n16899_o = 2'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b11;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b10;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b11;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16915_o = 2'b10;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16915_o = 2'b10;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16915_o = 2'b10;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16915_o = 2'b10;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16915_o = 2'b11;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16915_o = 2'b01;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16915_o = 2'b11;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16915_o = 2'b10;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16915_o = 2'b10;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16915_o = n16101_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16915_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16915_o = 2'b00;
      default: n16915_o = 2'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b10;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b10;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16925_o = 2'b01;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16925_o = 2'b10;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16925_o = 2'b01;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16925_o = 2'b11;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16925_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16925_o = 2'b00;
      default: n16925_o = 2'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b1;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b1;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16934_o = 1'b1;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16934_o = 1'b1;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16934_o = 1'b1;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16934_o = n16004_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16934_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16934_o = 1'b0;
      default: n16934_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n13151_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16937_o = 7'b1001111;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n13151_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n16697_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n16666_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n16628_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n16549_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n16504_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n16482_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n16467_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16937_o = 7'b1000100;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n13151_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n13151_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16937_o = n16387_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16937_o = 7'b0111101;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16937_o = n16349_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16937_o = 7'b0111011;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16937_o = 7'b1000000;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16937_o = n16279_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16937_o = 7'b0111000;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16937_o = n16264_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16937_o = n16257_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16937_o = n16248_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16937_o = n16226_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16937_o = 7'b0110011;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16937_o = n16214_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16937_o = n16207_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16937_o = 7'b0110000;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16937_o = 7'b0101111;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16937_o = 7'b1000001;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16937_o = n16176_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16937_o = 7'b1000001;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16937_o = 7'b1000000;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16937_o = n16144_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16937_o = n16137_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16937_o = n16125_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16937_o = n16111_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16937_o = n16093_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16937_o = n16069_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16937_o = 7'b0100100;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16937_o = n16007_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16937_o = 7'b0100010;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16937_o = 7'b0100001;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16937_o = n15989_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16937_o = n15971_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16937_o = 7'b0000000;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16937_o = 7'b0011101;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16937_o = n15923_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16937_o = 7'b0011011;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16937_o = 7'b0011010;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16937_o = 7'b0011001;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16937_o = n15822_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16937_o = 7'b1001101;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16937_o = 7'b0100101;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16937_o = 7'b1001011;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16937_o = n15777_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16937_o = 7'b1001001;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16937_o = n15699_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16937_o = n15418_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16937_o = n15349_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16937_o = n15300_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16937_o = 7'b1001111;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16937_o = n15213_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16937_o = n15083_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16937_o = n14951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16937_o = n14804_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16937_o = n14771_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16937_o = n14691_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16937_o = n14638_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16937_o = 7'b0000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16937_o = 7'b0000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16937_o = 7'b0000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16937_o = 7'b0000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16937_o = 7'b0000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16937_o = 7'b0000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16937_o = n14160_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16937_o = 7'b0000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16937_o = n13911_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16937_o = 7'b0000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16937_o = n13736_o;
      default: n16937_o = 7'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16939_o = n16177_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16939_o = 1'b1;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16939_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16939_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16939_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16939_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16939_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16939_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16939_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16939_o = n14161_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16939_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16939_o = n13912_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16939_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16939_o = 1'b0;
      default: n16939_o = 1'bX;
    endcase
  assign n16940_o = n13837_o[0];
  assign n16941_o = n14466_o[0];
  assign n16942_o = n14506_o[0];
  assign n16943_o = n14532_o[0];
  assign n16944_o = r[127];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16946_o = n16943_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16946_o = n16942_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16946_o = n16941_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16946_o = n14345_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16946_o = n16944_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16946_o = n16940_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16946_o = n16944_o;
      default: n16946_o = 1'bX;
    endcase
  assign n16947_o = n13837_o[1];
  assign n16948_o = n14466_o[1];
  assign n16949_o = n14506_o[1];
  assign n16950_o = n14532_o[1];
  assign n16951_o = r[128];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16953_o = n16950_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16953_o = n16949_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16953_o = n16948_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16953_o = n14340_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16953_o = n16951_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16953_o = n16947_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16953_o = n16951_o;
      default: n16953_o = 1'bX;
    endcase
  assign n16954_o = n13837_o[2];
  assign n16955_o = n14466_o[2];
  assign n16956_o = n14532_o[2];
  assign n16957_o = r[129];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16959_o = n16956_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16959_o = n16955_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16959_o = n14335_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16959_o = n16957_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16959_o = n16954_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16959_o = n16957_o;
      default: n16959_o = 1'bX;
    endcase
  assign n16960_o = n13837_o[3];
  assign n16961_o = n14466_o[3];
  assign n16962_o = n14508_o[0];
  assign n16963_o = n14532_o[3];
  assign n16964_o = r[130];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16966_o = n16963_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16966_o = n16962_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16966_o = n16961_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16966_o = n14330_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16966_o = n16964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16966_o = n16960_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16966_o = n16964_o;
      default: n16966_o = 1'bX;
    endcase
  assign n16967_o = n13837_o[4];
  assign n16968_o = n14466_o[4];
  assign n16969_o = n14508_o[1];
  assign n16970_o = n14536_o[0];
  assign n16971_o = r[131];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16973_o = n16970_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16973_o = n16969_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16973_o = n16968_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16973_o = n14325_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16973_o = n16971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16973_o = n16967_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16973_o = n16971_o;
      default: n16973_o = 1'bX;
    endcase
  assign n16974_o = n13837_o[5];
  assign n16975_o = n14466_o[5];
  assign n16976_o = n14508_o[2];
  assign n16977_o = n14536_o[1];
  assign n16978_o = r[132];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16980_o = n16977_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16980_o = n16976_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16980_o = n16975_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16980_o = n14320_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16980_o = n16978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16980_o = n16974_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16980_o = n16978_o;
      default: n16980_o = 1'bX;
    endcase
  assign n16981_o = n13837_o[6];
  assign n16982_o = n14466_o[6];
  assign n16983_o = n14508_o[3];
  assign n16984_o = n14536_o[2];
  assign n16985_o = r[133];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16987_o = n16984_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16987_o = n16983_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16987_o = n16982_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16987_o = n14315_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16987_o = n16985_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16987_o = n16981_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16987_o = n16985_o;
      default: n16987_o = 1'bX;
    endcase
  assign n16988_o = n13837_o[7];
  assign n16989_o = n14466_o[7];
  assign n16990_o = n14508_o[4];
  assign n16991_o = n14536_o[3];
  assign n16992_o = r[134];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n16994_o = n16991_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n16994_o = n16990_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n16994_o = n16989_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n16994_o = n14310_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n16994_o = n16992_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n16994_o = n16988_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n16994_o = n16992_o;
      default: n16994_o = 1'bX;
    endcase
  assign n16995_o = n13837_o[8];
  assign n16996_o = n14466_o[8];
  assign n16997_o = n14540_o[0];
  assign n16998_o = r[135];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17000_o = 1'b1;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16424_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17000_o = n16997_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17000_o = n16996_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17000_o = n14305_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17000_o = n16998_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17000_o = n16995_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17000_o = n16998_o;
      default: n17000_o = 1'bX;
    endcase
  assign n17001_o = n13837_o[9];
  assign n17002_o = n14466_o[9];
  assign n17003_o = n14540_o[1];
  assign n17004_o = r[136];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17006_o = n15421_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17006_o = n15303_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17006_o = n17003_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17006_o = n17002_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17006_o = n14300_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17006_o = n17004_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17006_o = n17001_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17006_o = n17004_o;
      default: n17006_o = 1'bX;
    endcase
  assign n17007_o = n13837_o[10];
  assign n17008_o = n14466_o[10];
  assign n17009_o = n14540_o[2];
  assign n17010_o = r[137];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17012_o = n17009_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17012_o = n17008_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17012_o = n14295_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17012_o = n17010_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17012_o = n17007_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17012_o = n17010_o;
      default: n17012_o = 1'bX;
    endcase
  assign n17013_o = n13837_o[11];
  assign n17014_o = n14466_o[11];
  assign n17015_o = n14540_o[3];
  assign n17016_o = r[138];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17018_o = n17015_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17018_o = n17014_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17018_o = n14290_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17018_o = n17016_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17018_o = n17013_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17018_o = n17016_o;
      default: n17018_o = 1'bX;
    endcase
  assign n17019_o = n13837_o[12];
  assign n17020_o = n14174_o[0];
  assign n17021_o = n14466_o[12];
  assign n17022_o = n14544_o[0];
  assign n17023_o = n15963_o[0];
  assign n17024_o = r[139];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17026_o = n17023_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17026_o = n17022_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17026_o = n17021_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17026_o = n14285_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17026_o = n17020_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17026_o = n17024_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17026_o = n17019_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17026_o = n17024_o;
      default: n17026_o = 1'bX;
    endcase
  assign n17027_o = n13837_o[13];
  assign n17028_o = n14174_o[1];
  assign n17029_o = n14466_o[13];
  assign n17030_o = n14544_o[1];
  assign n17031_o = n15963_o[1];
  assign n17032_o = r[140];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17034_o = n17031_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17034_o = n17030_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17034_o = n17029_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17034_o = n14280_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17034_o = n17028_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17034_o = n17032_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17034_o = n17027_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17034_o = n17032_o;
      default: n17034_o = 1'bX;
    endcase
  assign n17035_o = n13837_o[14];
  assign n17036_o = n14174_o[2];
  assign n17037_o = n14466_o[14];
  assign n17038_o = n14544_o[2];
  assign n17039_o = n15963_o[2];
  assign n17040_o = r[141];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17042_o = n17039_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17042_o = n17038_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17042_o = n17037_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17042_o = n14275_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17042_o = n17036_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17042_o = n17040_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17042_o = n17035_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17042_o = n17040_o;
      default: n17042_o = 1'bX;
    endcase
  assign n17043_o = n13837_o[15];
  assign n17044_o = n14174_o[3];
  assign n17045_o = n14466_o[15];
  assign n17046_o = n14544_o[3];
  assign n17047_o = n15963_o[3];
  assign n17048_o = r[142];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17050_o = n17047_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17050_o = n17046_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17050_o = n17045_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17050_o = n14270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17050_o = n17044_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17050_o = n17048_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17050_o = n17043_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17050_o = n17048_o;
      default: n17050_o = 1'bX;
    endcase
  assign n17051_o = n13837_o[16];
  assign n17052_o = n14466_o[16];
  assign n17053_o = n14548_o[0];
  assign n17054_o = r[143];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17056_o = n17053_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17056_o = n17052_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17056_o = n14265_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17056_o = n17054_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17056_o = n17051_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17056_o = n17054_o;
      default: n17056_o = 1'bX;
    endcase
  assign n17057_o = n13837_o[17];
  assign n17058_o = n14466_o[17];
  assign n17059_o = n14548_o[1];
  assign n17060_o = n16336_o[0];
  assign n17061_o = n16551_o[0];
  assign n17062_o = n16611_o[0];
  assign n17063_o = r[144];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17062_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17061_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17060_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17065_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17065_o = n17059_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17065_o = n17058_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17065_o = n14260_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17065_o = n17063_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17065_o = n17057_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17065_o = n17063_o;
      default: n17065_o = 1'bX;
    endcase
  assign n17066_o = n13837_o[18];
  assign n17067_o = n14466_o[18];
  assign n17068_o = n14548_o[2];
  assign n17069_o = n16336_o[1];
  assign n17070_o = n16551_o[1];
  assign n17071_o = n16611_o[1];
  assign n17072_o = r[145];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17071_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17070_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17069_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17074_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17074_o = n17068_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17074_o = n17067_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17074_o = n14255_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17074_o = n17072_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17074_o = n17066_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17074_o = n17072_o;
      default: n17074_o = 1'bX;
    endcase
  assign n17075_o = n13837_o[19];
  assign n17076_o = n14466_o[19];
  assign n17077_o = n14548_o[3];
  assign n17078_o = r[146];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17080_o = n17077_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17080_o = n17076_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17080_o = n14250_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17080_o = n14162_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17080_o = n17078_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17080_o = n17075_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17080_o = n17078_o;
      default: n17080_o = 1'bX;
    endcase
  assign n17081_o = n13837_o[20];
  assign n17082_o = n14466_o[20];
  assign n17083_o = n14552_o[0];
  assign n17084_o = r[147];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17086_o = n15701_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17086_o = n15085_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17086_o = n17083_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17086_o = n17082_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17086_o = n14245_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17086_o = n17084_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17086_o = n17081_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17086_o = n17084_o;
      default: n17086_o = 1'bX;
    endcase
  assign n17087_o = n13837_o[21];
  assign n17088_o = n14466_o[21];
  assign n17089_o = n14552_o[1];
  assign n17090_o = n15215_o[0];
  assign n17091_o = r[148];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17093_o = n17090_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17093_o = n17089_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17093_o = n17088_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17093_o = n14240_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17093_o = n17091_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17093_o = n17087_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17093_o = n17091_o;
      default: n17093_o = 1'bX;
    endcase
  assign n17094_o = n13837_o[22];
  assign n17095_o = n14466_o[22];
  assign n17096_o = n14552_o[2];
  assign n17097_o = n15215_o[1];
  assign n17098_o = r[149];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17100_o = n17097_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17100_o = n17096_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17100_o = n17095_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17100_o = n14235_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17100_o = n17098_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17100_o = n17094_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17100_o = n17098_o;
      default: n17100_o = 1'bX;
    endcase
  assign n17101_o = n13837_o[23];
  assign n17102_o = n14466_o[23];
  assign n17103_o = n14552_o[3];
  assign n17104_o = r[150];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17106_o = n15703_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17106_o = n14953_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17106_o = n17103_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17106_o = n17102_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17106_o = n14230_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17106_o = n17104_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17106_o = n17101_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17106_o = n17104_o;
      default: n17106_o = 1'bX;
    endcase
  assign n17107_o = n13837_o[24];
  assign n17108_o = n14466_o[24];
  assign n17109_o = n14556_o[0];
  assign n17110_o = r[151];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n16742_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17112_o = n14715_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17112_o = n14665_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17112_o = n14609_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17112_o = n17109_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17112_o = n17108_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17112_o = n14225_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17112_o = n14164_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17112_o = n17110_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17112_o = n17107_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17112_o = n17110_o;
      default: n17112_o = 1'bX;
    endcase
  assign n17113_o = n13837_o[25];
  assign n17114_o = n14466_o[25];
  assign n17115_o = n14556_o[1];
  assign n17116_o = r[152];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n16641_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n16553_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n16426_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17118_o = n16389_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17118_o = n17115_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17118_o = n17114_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17118_o = n14220_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17118_o = n17116_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17118_o = n17113_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17118_o = n17116_o;
      default: n17118_o = 1'bX;
    endcase
  assign n17119_o = n13837_o[26];
  assign n17120_o = n14466_o[26];
  assign n17121_o = n14556_o[2];
  assign n17122_o = r[153];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17124_o = n17121_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17124_o = n17120_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17124_o = n14215_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17124_o = n17122_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17124_o = n17119_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17124_o = n17122_o;
      default: n17124_o = 1'bX;
    endcase
  assign n17125_o = n13837_o[27];
  assign n17126_o = n14466_o[27];
  assign n17127_o = n14556_o[3];
  assign n17128_o = r[154];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n16639_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n16506_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17130_o = n17127_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17130_o = n17126_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17130_o = n14210_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17130_o = n17128_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17130_o = n17125_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17130_o = n17128_o;
      default: n17130_o = 1'bX;
    endcase
  assign n17131_o = n13837_o[28];
  assign n17132_o = n14466_o[28];
  assign n17133_o = n14560_o[0];
  assign n17134_o = r[155];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17136_o = 1'b1;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17136_o = n17133_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17136_o = n17132_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17136_o = n14205_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17136_o = n17134_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17136_o = n17131_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17136_o = n17134_o;
      default: n17136_o = 1'bX;
    endcase
  assign n17137_o = n13837_o[29];
  assign n17138_o = n14466_o[29];
  assign n17139_o = n14560_o[1];
  assign n17140_o = r[156];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17142_o = n17139_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17142_o = n17138_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17142_o = n14200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17142_o = n17140_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17142_o = n17137_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17142_o = n17140_o;
      default: n17142_o = 1'bX;
    endcase
  assign n17143_o = n13837_o[30];
  assign n17144_o = n14466_o[30];
  assign n17145_o = n14560_o[2];
  assign n17146_o = r[157];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17148_o = n17145_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17148_o = n17144_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17148_o = n14195_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17148_o = n17146_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17148_o = n17143_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17148_o = n17146_o;
      default: n17148_o = 1'bX;
    endcase
  assign n17149_o = n13837_o[31];
  assign n17150_o = n14466_o[31];
  assign n17151_o = n14560_o[3];
  assign n17152_o = r[158];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17154_o = n17151_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17154_o = n17150_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17154_o = n14190_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17154_o = n17152_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17154_o = n17149_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17154_o = n17152_o;
      default: n17154_o = 1'bX;
    endcase
  assign n17155_o = r[519];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17157_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n16455_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17157_o = n16288_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17157_o = n16153_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17157_o = s_nz;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17157_o = n17155_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17157_o = 1'b0;
      default: n17157_o = 1'bX;
    endcase
  assign n17158_o = n16051_o[0];
  assign n17159_o = n16699_o[0];
  assign n17160_o = r[648];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n16803_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17159_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17162_o = n17158_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17162_o = n16025_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17162_o = n15980_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17162_o = n15925_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17162_o = n15705_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17162_o = n15369_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17162_o = n15322_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17162_o = n15251_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17162_o = n15107_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17162_o = n14978_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17162_o = n14954_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17162_o = n14793_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17162_o = n14701_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17162_o = n14651_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17162_o = n14595_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17162_o = n14586_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17162_o = n17160_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17162_o = n17160_o;
      default: n17162_o = 1'bX;
    endcase
  assign n17163_o = n16051_o[2:1];
  assign n17164_o = n16699_o[2:1];
  assign n17165_o = r[650:649];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n16804_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17164_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n16556_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17167_o = n17163_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17167_o = n15928_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17167_o = n15707_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17167_o = n15423_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17167_o = n15351_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17167_o = n15249_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17167_o = n15216_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17167_o = n14980_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17167_o = n14813_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17167_o = n14795_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17167_o = n14699_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17167_o = n14649_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17167_o = n14593_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17167_o = n14566_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17167_o = n17165_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17167_o = n17165_o;
      default: n17167_o = 2'bX;
    endcase
  assign n17168_o = n15709_o[12:0];
  assign n17169_o = r[663:651];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n16805_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n16558_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n16508_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17171_o = n16269_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17171_o = n16185_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17171_o = n15837_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17171_o = n13526_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17171_o = n15795_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17171_o = n13526_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17171_o = n17168_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17171_o = n15426_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17171_o = n15354_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17171_o = n15306_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17171_o = n15112_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17171_o = n15087_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17171_o = n14815_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17171_o = 13'b0000000110110;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17171_o = n14703_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17171_o = n14653_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17171_o = n14597_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17171_o = n14568_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17171_o = n13976_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17171_o = n17169_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17171_o = n17169_o;
      default: n17171_o = 13'bX;
    endcase
  assign n17172_o = n15709_o[25:13];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17174_o = n16700_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17174_o = n16629_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17174_o = n16483_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17174_o = n16468_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b1111111111110;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000001;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17174_o = 13'b1111111111111;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000001;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17174_o = n16178_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000001;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17174_o = 13'b0000000111000;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17174_o = n15995_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17174_o = n15984_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17174_o = 13'b1111111111111;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17174_o = n15835_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17174_o = n17172_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17174_o = 13'b0000000000001;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17174_o = n15308_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17174_o = n14863_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17174_o = n14773_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17174_o = n14690_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17174_o = n14639_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17174_o = 13'b0000000000000;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17174_o = 13'b0000000000000;
      default: n17174_o = 13'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17176_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17176_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17176_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17176_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17176_o = 1'b0;
      default: n17176_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17178_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17178_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17178_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17178_o = n13471_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17178_o = n13471_o;
      default: n17178_o = 1'bX;
    endcase
  assign n17179_o = n13828_o[0];
  assign n17180_o = n14165_o[0];
  assign n17181_o = n15961_o[0];
  assign n17182_o = r[679];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17184_o = n17181_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17184_o = n17182_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17184_o = n17180_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17184_o = n13970_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17184_o = n13917_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17184_o = n17179_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17184_o = n17182_o;
      default: n17184_o = 1'bX;
    endcase
  assign n17185_o = n13828_o[1];
  assign n17186_o = n14165_o[1];
  assign n17187_o = n15961_o[1];
  assign n17188_o = r[680];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17190_o = n16161_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17190_o = n17187_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17190_o = n17188_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17190_o = n17186_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17190_o = n13969_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17190_o = n13914_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17190_o = n17185_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17190_o = n17188_o;
      default: n17190_o = 1'bX;
    endcase
  assign n17191_o = n13828_o[2];
  assign n17192_o = n14165_o[2];
  assign n17193_o = n15961_o[2];
  assign n17194_o = r[681];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17196_o = n17193_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17196_o = n17194_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17196_o = n17192_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17196_o = n13942_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17196_o = n13869_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17196_o = n17191_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17196_o = n17194_o;
      default: n17196_o = 1'bX;
    endcase
  assign n17197_o = n13828_o[3];
  assign n17198_o = n14165_o[3];
  assign n17199_o = n15961_o[3];
  assign n17200_o = r[682];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17202_o = n17199_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17202_o = n17200_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17202_o = n17198_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17202_o = n13943_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17202_o = n13870_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17202_o = n17197_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17202_o = n17200_o;
      default: n17202_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17204_o = n13558_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17204_o = n13749_o;
      default: n17204_o = 5'bX;
    endcase
  assign n17205_o = n13465_o[0];
  assign n17206_o = r[697];
  /* fpu.vhdl:650:9  */
  assign n17207_o = n13152_o ? n17205_o : n17206_o;
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17209_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17209_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17209_o = n17207_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17209_o = n17207_o;
      default: n17209_o = 1'bX;
    endcase
  assign n17210_o = n13465_o[1];
  assign n17211_o = r[698];
  /* fpu.vhdl:650:9  */
  assign n17212_o = n13152_o ? n17210_o : n17211_o;
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17214_o = 1'b1;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17214_o = n17212_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17214_o = n17212_o;
      default: n17214_o = 1'bX;
    endcase
  assign n17215_o = n13465_o[2];
  assign n17216_o = r[699];
  /* fpu.vhdl:650:9  */
  assign n17217_o = n13152_o ? n17215_o : n17216_o;
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n16704_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17219_o = n17217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17219_o = n17217_o;
      default: n17219_o = 1'bX;
    endcase
  assign n17220_o = n13465_o[5:3];
  assign n17221_o = r[702:700];
  /* fpu.vhdl:650:9  */
  assign n17222_o = n13152_o ? n17220_o : n17221_o;
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17224_o = n14643_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17224_o = n17222_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17224_o = n13740_o;
      default: n17224_o = 3'bX;
    endcase
  assign n17225_o = n13465_o[6];
  assign n17226_o = r[703];
  /* fpu.vhdl:650:9  */
  assign n17227_o = n13152_o ? n17225_o : n17226_o;
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17229_o = n15713_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17229_o = n14959_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17229_o = n17227_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17229_o = n17227_o;
      default: n17229_o = 1'bX;
    endcase
  assign n17230_o = n13465_o[8];
  assign n17231_o = r[705];
  /* fpu.vhdl:650:9  */
  assign n17232_o = n13152_o ? n17230_o : n17231_o;
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17234_o = n15826_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17234_o = n15781_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17234_o = n17232_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17234_o = n17232_o;
      default: n17234_o = 1'bX;
    endcase
  assign n17235_o = n13465_o[9];
  assign n17236_o = r[706];
  /* fpu.vhdl:650:9  */
  assign n17237_o = n13152_o ? n17235_o : n17236_o;
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17239_o = n14963_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17239_o = n17237_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17239_o = n17237_o;
      default: n17239_o = 1'bX;
    endcase
  assign n17240_o = n13744_o[0];
  assign n17241_o = n13465_o[10];
  assign n17242_o = r[707];
  /* fpu.vhdl:650:9  */
  assign n17243_o = n13152_o ? n17241_o : n17242_o;
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17245_o = n15717_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17245_o = n17243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17245_o = n17240_o;
      default: n17245_o = 1'bX;
    endcase
  assign n17246_o = n13744_o[1];
  assign n17247_o = n13465_o[11];
  assign n17248_o = r[708];
  /* fpu.vhdl:650:9  */
  assign n17249_o = n13152_o ? n17247_o : n17248_o;
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17251_o = n17249_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17251_o = n17246_o;
      default: n17251_o = 1'bX;
    endcase
  assign n17252_o = n16113_o[0];
  assign n17253_o = n16250_o[0];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b1;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17255_o = n16258_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17255_o = n17253_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17255_o = n16227_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17255_o = 1'b1;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17255_o = n16208_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17255_o = 1'b1;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17255_o = n16138_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17255_o = n16126_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17255_o = n17252_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17255_o = 1'b1;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17255_o = 1'b1;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17255_o = n15827_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17255_o = n15782_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17255_o = n15217_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17255_o = n13915_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17255_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17255_o = 1'b0;
      default: n17255_o = 1'bX;
    endcase
  assign n17256_o = n16113_o[2:1];
  assign n17257_o = n16250_o[2:1];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17259_o = n17257_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17259_o = 2'b00;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17259_o = n17256_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17259_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17259_o = n13562_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17259_o = n13562_o;
      default: n17259_o = 2'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17261_o = n16179_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17261_o = n13916_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17261_o = n13477_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17261_o = n13477_o;
      default: n17261_o = 2'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17263_o = n16769_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17263_o = n15846_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17263_o = n15828_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17263_o = 2'b10;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17263_o = n15770_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17263_o = n15732_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17263_o = n15718_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17263_o = n15243_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17263_o = n15088_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17263_o = n14964_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17263_o = n14166_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17263_o = 2'b00;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17263_o = n13745_o;
      default: n17263_o = 2'bX;
    endcase
  assign n17264_o = r[716];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17266_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17266_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17266_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17266_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17266_o = n17264_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17266_o = 1'b0;
      default: n17266_o = 1'bX;
    endcase
  assign n17267_o = r[717];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17269_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17269_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17269_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17269_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17269_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17269_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17269_o = n17267_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17269_o = 1'b0;
      default: n17269_o = 1'bX;
    endcase
  assign n17270_o = r[718];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17272_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17272_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17272_o = n17270_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17272_o = 1'b0;
      default: n17272_o = 1'bX;
    endcase
  assign n17273_o = r[719];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17275_o = n17273_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17275_o = 1'b0;
      default: n17275_o = 1'bX;
    endcase
  assign n17276_o = r[720];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17278_o = n15720_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17278_o = n15090_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17278_o = n14966_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17278_o = n17276_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17278_o = 1'b0;
      default: n17278_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17280_o = n15990_o;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17280_o = n15842_o;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17280_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17280_o = n14864_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17280_o = n13479_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17280_o = n13479_o;
      default: n17280_o = 1'bX;
    endcase
  assign n17313_o = r[518:399];
  assign n17315_o = r[647:520];
  assign n17338_o = n13465_o[7];
  assign n17339_o = r[704];
  /* fpu.vhdl:650:9  */
  assign n17340_o = n13152_o ? n17338_o : n17339_o;
  assign n17351_o = n14514_o[3:0];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17354_o = n17351_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17354_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17354_o = n13830_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17354_o = 4'b1111;
      default: n17354_o = 4'bX;
    endcase
  assign n17355_o = n14514_o[7:4];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17358_o = n17355_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17358_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17358_o = n13821_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17358_o = 4'b1111;
      default: n17358_o = 4'bX;
    endcase
  assign n17359_o = n14514_o[11:8];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17362_o = n17359_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17362_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17362_o = n13812_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17362_o = 4'b1111;
      default: n17362_o = 4'bX;
    endcase
  assign n17363_o = n14514_o[15:12];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17366_o = n17363_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17366_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17366_o = n13803_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17366_o = 4'b1111;
      default: n17366_o = 4'bX;
    endcase
  assign n17367_o = n14514_o[19:16];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17370_o = n17367_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17370_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17370_o = n13794_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17370_o = 4'b1111;
      default: n17370_o = 4'bX;
    endcase
  assign n17371_o = n14514_o[23:20];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17374_o = n17371_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17374_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17374_o = n13785_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17374_o = 4'b1111;
      default: n17374_o = 4'bX;
    endcase
  assign n17375_o = n14514_o[27:24];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17378_o = n17375_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17378_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17378_o = n13776_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17378_o = 4'b1111;
      default: n17378_o = 4'bX;
    endcase
  assign n17379_o = n14514_o[31:28];
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17382_o = n17379_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17382_o = 4'b1111;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17382_o = n13767_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17382_o = 4'b1111;
      default: n17382_o = 4'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17393_o = n14517_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17393_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17393_o = n13747_o;
      default: n17393_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17407_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17407_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17407_o = 1'b0;
      default: n17407_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b1;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b1;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17415_o = n16706_o;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17415_o = n16667_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17415_o = n16631_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17415_o = n16561_o;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b1;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b1;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17415_o = n16392_o;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17415_o = n16073_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17415_o = n15930_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17415_o = n15722_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17415_o = n15431_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17415_o = n15359_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17415_o = n15313_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17415_o = n15219_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17415_o = n15092_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17415_o = n14969_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17415_o = n14807_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17415_o = n14777_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17415_o = n14695_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17415_o = n14645_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17415_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17415_o = 1'b0;
      default: n17415_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17420_o = n16745_o;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b1;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17420_o = n16429_o;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17420_o = n14718_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17420_o = n14668_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17420_o = n14612_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17420_o = n14168_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17420_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17420_o = 1'b0;
      default: n17420_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17424_o = n15435_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17424_o = n15363_o;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17424_o = n15221_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17424_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17424_o = 1'b0;
      default: n17424_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17433_o = n16669_o;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17433_o = n16633_o;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17433_o = n16510_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17433_o = n16471_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17433_o = n16075_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17433_o = n15932_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17433_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17433_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17433_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17433_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17433_o = 1'b0;
      default: n17433_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17442_o = n16513_o;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b1;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17442_o = n16474_o;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b1;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b1;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17442_o = n15934_o;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17442_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17442_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17442_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17442_o = 1'b0;
      default: n17442_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17454_o = 1'b1;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17454_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17454_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17454_o = 1'b0;
      default: n17454_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17459_o = n16276_o;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17459_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17459_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17459_o = 1'b0;
      default: n17459_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17464_o = 1'b1;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17464_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17464_o = 1'b0;
      default: n17464_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17468_o = n16230_o;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17468_o = n16200_o;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17468_o = n16129_o;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17468_o = n16102_o;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17468_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17468_o = 1'b0;
      default: n17468_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17476_o = n16077_o;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17476_o = n16028_o;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17476_o = 1'b1;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17476_o = 1'b1;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17476_o = 1'b1;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17476_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17476_o = 1'b1;
      default: n17476_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17480_o = n15724_o;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17480_o = n15438_o;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17480_o = n15316_o;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17480_o = n15223_o;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17480_o = n15094_o;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17480_o = n14971_o;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17480_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17480_o = 1'b0;
      default: n17480_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b1;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b1;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17493_o = 1'b1;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17493_o = 1'b1;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17493_o = 1'b1;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17493_o = 1'b1;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17493_o = 1'b1;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17493_o = 1'b1;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17493_o = 1'b1;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17493_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17493_o = 1'b0;
      default: n17493_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17497_o = n15786_o;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17497_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17497_o = 1'b0;
      default: n17497_o = 1'bX;
    endcase
  /* fpu.vhdl:776:9  */
  always @*
    case (n16808_o)
      80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b1;
      80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010: n17504_o = 1'b0;
      80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001: n17504_o = 1'b0;
      default: n17504_o = 1'bX;
    endcase
  /* fpu.vhdl:2286:9  */
  assign n17509_o = n17424_o ? 1'b1 : n17124_o;
  /* fpu.vhdl:2289:9  */
  assign n17513_o = n17480_o ? 2'b11 : n16836_o;
  assign n17515_o = {n16881_o, n16872_o};
  /* fpu.vhdl:2289:9  */
  assign n17516_o = n17480_o ? 4'b0001 : n17515_o;
  assign n17517_o = {2'b11, 1'b0};
  assign n17518_o = {n17167_o, n17162_o};
  /* fpu.vhdl:2289:9  */
  assign n17519_o = n17480_o ? n17517_o : n17518_o;
  /* fpu.vhdl:2289:9  */
  assign n17521_o = n17480_o ? 1'b1 : n17415_o;
  /* fpu.vhdl:2289:9  */
  assign n17523_o = n17480_o ? 1'b1 : n17420_o;
  /* fpu.vhdl:2297:9  */
  assign n17525_o = n17523_o ? 1'b1 : n17275_o;
  assign n17526_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, 1'b0, n17204_o, n13473_o, n17202_o, n17196_o, n17190_o, n17184_o, n17178_o, n17176_o, n17174_o, n17171_o, n17519_o, n17315_o, n17157_o, n17313_o, n13469_o, n17154_o, n17148_o, n17142_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n17056_o, n17050_o, n17042_o, n17034_o, n17026_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n13556_o, n16939_o, 1'b0, n16937_o};
  /* fpu.vhdl:2303:19  */
  assign n17527_o = n17526_o[719];
  /* fpu.vhdl:2303:38  */
  assign n17528_o = r[134];
  /* fpu.vhdl:2303:27  */
  assign n17529_o = n17527_o & n17528_o;
  /* fpu.vhdl:2303:50  */
  assign n17530_o = ~n17529_o;
  /* fpu.vhdl:2304:41  */
  assign n17531_o = r[131];
  /* fpu.vhdl:2304:30  */
  assign n17532_o = n17424_o & n17531_o;
  /* fpu.vhdl:2304:53  */
  assign n17533_o = ~n17532_o;
  /* fpu.vhdl:2303:56  */
  assign n17534_o = n17530_o & n17533_o;
  /* fpu.vhdl:2300:9  */
  assign n17537_o = n17543_o ? 1'b1 : n17176_o;
  /* fpu.vhdl:2300:9  */
  assign n17538_o = n17544_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:2300:9  */
  assign n17541_o = n17521_o ? 7'b0000000 : n16937_o;
  /* fpu.vhdl:2300:9  */
  assign n17542_o = n17521_o ? 1'b1 : n16939_o;
  /* fpu.vhdl:2300:9  */
  assign n17543_o = n17521_o & n17534_o;
  /* fpu.vhdl:2300:9  */
  assign n17544_o = n17521_o & n17534_o;
  /* fpu.vhdl:2300:9  */
  assign n17546_o = n17521_o ? 1'b1 : n17407_o;
  /* fpu.vhdl:2316:52  */
  assign n17547_o = r[236:175];
  /* fpu.vhdl:2316:66  */
  assign n17549_o = {n17547_o, 2'b00};
  /* fpu.vhdl:2315:13  */
  assign n17551_o = msel_1 == 2'b00;
  /* fpu.vhdl:2318:52  */
  assign n17552_o = r[316:255];
  /* fpu.vhdl:2318:66  */
  assign n17554_o = {n17552_o, 2'b00};
  /* fpu.vhdl:2317:13  */
  assign n17556_o = msel_1 == 2'b01;
  /* fpu.vhdl:2320:42  */
  assign n17557_o = r[647:584];
  /* fpu.vhdl:2319:13  */
  assign n17559_o = msel_1 == 2'b10;
  /* fpu.vhdl:2322:43  */
  assign n17560_o = r[460:399];
  /* fpu.vhdl:2322:57  */
  assign n17562_o = {n17560_o, 2'b00};
  assign n17563_o = {n17559_o, n17556_o, n17551_o};
  /* fpu.vhdl:2314:9  */
  always @*
    case (n17563_o)
      3'b100: n17564_o = n17557_o;
      3'b010: n17564_o = n17554_o;
      3'b001: n17564_o = n17549_o;
      default: n17564_o = n17562_o;
    endcase
  /* fpu.vhdl:2326:52  */
  assign n17565_o = r[396:335];
  /* fpu.vhdl:2326:66  */
  assign n17567_o = {n17565_o, 2'b00};
  /* fpu.vhdl:2325:13  */
  assign n17569_o = msel_2 == 2'b00;
  /* fpu.vhdl:2328:46  */
  assign n17571_o = {8'b00000000, inverse_est};
  /* fpu.vhdl:2328:60  */
  assign n17573_o = {n17571_o, 1'b0};
  /* fpu.vhdl:2328:66  */
  assign n17575_o = {n17573_o, 36'b000000000000000000000000000000000000};
  /* fpu.vhdl:2327:13  */
  assign n17577_o = msel_2 == 2'b01;
  /* fpu.vhdl:2330:42  */
  assign n17578_o = r[583:520];
  /* fpu.vhdl:2329:13  */
  assign n17580_o = msel_2 == 2'b10;
  /* fpu.vhdl:2332:43  */
  assign n17581_o = r[460:399];
  /* fpu.vhdl:2332:57  */
  assign n17583_o = {n17581_o, 2'b00};
  assign n17584_o = {n17580_o, n17577_o, n17569_o};
  /* fpu.vhdl:2324:9  */
  always @*
    case (n17584_o)
      3'b100: n17585_o = n17578_o;
      3'b010: n17585_o = n17575_o;
      3'b001: n17585_o = n17567_o;
      default: n17585_o = n17583_o;
    endcase
  /* fpu.vhdl:2338:22  */
  assign n17586_o = r[708];
  /* fpu.vhdl:2338:30  */
  assign n17587_o = ~n17586_o;
  /* fpu.vhdl:2338:17  */
  assign n17591_o = n17587_o ? 2'b00 : 2'b11;
  /* fpu.vhdl:2338:17  */
  assign n17593_o = n17587_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:2336:13  */
  assign n17595_o = msel_add == 2'b01;
  /* fpu.vhdl:2345:45  */
  assign n17596_o = r[238:159];
  /* fpu.vhdl:2345:47  */
  assign n17597_o = n17596_o[79:16];
  /* fpu.vhdl:2343:13  */
  assign n17599_o = msel_add == 2'b10;
  /* fpu.vhdl:2348:41  */
  assign n17600_o = r[462:399];
  /* fpu.vhdl:2348:37  */
  assign n17602_o = {6'b000000, n17600_o};
  /* fpu.vhdl:2348:47  */
  assign n17603_o = r[518:463];
  /* fpu.vhdl:2348:43  */
  assign n17604_o = {n17602_o, n17603_o};
  /* fpu.vhdl:2348:49  */
  assign n17606_o = {n17604_o, 2'b00};
  /* fpu.vhdl:2346:13  */
  assign n17608_o = msel_add == 2'b11;
  assign n17609_o = {n17608_o, n17599_o, n17595_o};
  assign n17610_o = n17606_o[57:0];
  /* fpu.vhdl:2335:9  */
  always @*
    case (n17609_o)
      3'b100: n17612_o = n17610_o;
      3'b010: n17612_o = 58'b0000000000000000000000000000000000000000000000000000000000;
      3'b001: n17612_o = 58'b0000000000000000000000000000000000000000000000000000000000;
      default: n17612_o = 58'b0000000000000000000000000000000000000000000000000000000000;
    endcase
  assign n17613_o = n17597_o[52:0];
  assign n17614_o = n17606_o[110:58];
  /* fpu.vhdl:2335:9  */
  always @*
    case (n17609_o)
      3'b100: n17616_o = n17614_o;
      3'b010: n17616_o = n17613_o;
      3'b001: n17616_o = 53'b00000000000000000000000000000000000000000000000000000;
      default: n17616_o = 53'b00000000000000000000000000000000000000000000000000000;
    endcase
  assign n17617_o = n17597_o[54:53];
  assign n17618_o = n17606_o[112:111];
  /* fpu.vhdl:2335:9  */
  always @*
    case (n17609_o)
      3'b100: n17620_o = n17618_o;
      3'b010: n17620_o = n17617_o;
      3'b001: n17620_o = n17591_o;
      default: n17620_o = 2'b00;
    endcase
  assign n17621_o = n17597_o[55];
  assign n17622_o = n17606_o[113];
  /* fpu.vhdl:2335:9  */
  always @*
    case (n17609_o)
      3'b100: n17624_o = n17622_o;
      3'b010: n17624_o = n17621_o;
      3'b001: n17624_o = n17593_o;
      default: n17624_o = 1'b0;
    endcase
  assign n17625_o = n17597_o[63:56];
  assign n17626_o = n17606_o[121:114];
  /* fpu.vhdl:2335:9  */
  always @*
    case (n17609_o)
      3'b100: n17628_o = n17626_o;
      3'b010: n17628_o = n17625_o;
      3'b001: n17628_o = 8'b00000000;
      default: n17628_o = 8'b00000000;
    endcase
  assign n17629_o = n17606_o[127:122];
  /* fpu.vhdl:2335:9  */
  always @*
    case (n17609_o)
      3'b100: n17631_o = n17629_o;
      3'b010: n17631_o = 6'b000000;
      3'b001: n17631_o = 6'b000000;
      default: n17631_o = 6'b000000;
    endcase
  assign n17638_o = {n17631_o, n17628_o, n17624_o, n17620_o, n17616_o, n17612_o};
  /* fpu.vhdl:2352:37  */
  assign n17639_o = ~n17638_o;
  assign n17640_o = {n17631_o, n17628_o, n17624_o, n17620_o, n17616_o, n17612_o};
  /* fpu.vhdl:2351:9  */
  assign n17641_o = msel_inv ? n17639_o : n17640_o;
  /* fpu.vhdl:2358:34  */
  assign n17642_o = f_to_multiply[128:65];
  assign n17643_o = r[647:584];
  /* fpu.vhdl:2357:9  */
  assign n17644_o = n17468_o ? n17642_o : n17643_o;
  assign n17645_o = r[583:520];
  /* fpu.vhdl:2360:26  */
  assign n17646_o = multiply_to_f[0];
  /* fpu.vhdl:2361:23  */
  assign n17647_o = ~n17493_o;
  /* fpu.vhdl:2362:44  */
  assign n17648_o = multiply_to_f[64:1];
  /* fpu.vhdl:2364:44  */
  assign n17649_o = multiply_to_f[120:57];
  /* fpu.vhdl:2361:13  */
  assign n17650_o = n17647_o ? n17648_o : n17649_o;
  /* fpu.vhdl:2360:9  */
  assign n17651_o = n17646_o ? n17650_o : n17645_o;
  /* fpu.vhdl:2371:14  */
  assign n17652_o = r[721];
  /* fpu.vhdl:2372:25  */
  assign n17653_o = r[676:664];
  /* fpu.vhdl:2372:31  */
  assign n17655_o = n17653_o + 13'b1111111100011;
  /* fpu.vhdl:2374:25  */
  assign n17656_o = r[676:664];
  /* fpu.vhdl:2371:9  */
  assign n17657_o = n17652_o ? n17655_o : n17656_o;
  /* fpu.vhdl:2376:19  */
  assign n17659_o = $signed(n17657_o) < $signed(13'b1111111000000);
  /* fpu.vhdl:2378:22  */
  assign n17661_o = $signed(n17657_o) >= $signed(13'b0000000000000);
  /* fpu.vhdl:2381:47  */
  assign n17663_o = n17657_o[5:0];
  /* fpu.vhdl:401:18  */
  assign n17670_o = $unsigned(6'b000000) >= $unsigned(n17663_o);
  /* fpu.vhdl:401:13  */
  assign n17673_o = n17670_o ? 1'b1 : 1'b0;
  /* fpu.vhdl:401:18  */
  assign n17677_o = $unsigned(6'b000001) >= $unsigned(n17663_o);
  assign n17679_o = n17674_o[62];
  /* fpu.vhdl:401:13  */
  assign n17680_o = n17677_o ? 1'b1 : n17679_o;
  /* fpu.vhdl:401:18  */
  assign n17683_o = $unsigned(6'b000010) >= $unsigned(n17663_o);
  assign n17685_o = n17674_o[61];
  /* fpu.vhdl:401:13  */
  assign n17686_o = n17683_o ? 1'b1 : n17685_o;
  /* fpu.vhdl:401:18  */
  assign n17689_o = $unsigned(6'b000011) >= $unsigned(n17663_o);
  assign n17691_o = n17674_o[60];
  /* fpu.vhdl:401:13  */
  assign n17692_o = n17689_o ? 1'b1 : n17691_o;
  /* fpu.vhdl:401:18  */
  assign n17695_o = $unsigned(6'b000100) >= $unsigned(n17663_o);
  assign n17697_o = n17674_o[59];
  /* fpu.vhdl:401:13  */
  assign n17698_o = n17695_o ? 1'b1 : n17697_o;
  /* fpu.vhdl:401:18  */
  assign n17701_o = $unsigned(6'b000101) >= $unsigned(n17663_o);
  assign n17703_o = n17674_o[58];
  /* fpu.vhdl:401:13  */
  assign n17704_o = n17701_o ? 1'b1 : n17703_o;
  /* fpu.vhdl:401:18  */
  assign n17707_o = $unsigned(6'b000110) >= $unsigned(n17663_o);
  assign n17709_o = n17674_o[57];
  /* fpu.vhdl:401:13  */
  assign n17710_o = n17707_o ? 1'b1 : n17709_o;
  /* fpu.vhdl:401:18  */
  assign n17713_o = $unsigned(6'b000111) >= $unsigned(n17663_o);
  assign n17715_o = n17674_o[56];
  /* fpu.vhdl:401:13  */
  assign n17716_o = n17713_o ? 1'b1 : n17715_o;
  /* fpu.vhdl:401:18  */
  assign n17719_o = $unsigned(6'b001000) >= $unsigned(n17663_o);
  assign n17721_o = n17674_o[55];
  /* fpu.vhdl:401:13  */
  assign n17722_o = n17719_o ? 1'b1 : n17721_o;
  /* fpu.vhdl:401:18  */
  assign n17725_o = $unsigned(6'b001001) >= $unsigned(n17663_o);
  assign n17727_o = n17674_o[54];
  /* fpu.vhdl:401:13  */
  assign n17728_o = n17725_o ? 1'b1 : n17727_o;
  /* fpu.vhdl:401:18  */
  assign n17731_o = $unsigned(6'b001010) >= $unsigned(n17663_o);
  assign n17733_o = n17674_o[53];
  /* fpu.vhdl:401:13  */
  assign n17734_o = n17731_o ? 1'b1 : n17733_o;
  /* fpu.vhdl:401:18  */
  assign n17737_o = $unsigned(6'b001011) >= $unsigned(n17663_o);
  assign n17739_o = n17674_o[52];
  /* fpu.vhdl:401:13  */
  assign n17740_o = n17737_o ? 1'b1 : n17739_o;
  /* fpu.vhdl:401:18  */
  assign n17743_o = $unsigned(6'b001100) >= $unsigned(n17663_o);
  assign n17745_o = n17674_o[51];
  /* fpu.vhdl:401:13  */
  assign n17746_o = n17743_o ? 1'b1 : n17745_o;
  /* fpu.vhdl:401:18  */
  assign n17749_o = $unsigned(6'b001101) >= $unsigned(n17663_o);
  assign n17751_o = n17674_o[50];
  /* fpu.vhdl:401:13  */
  assign n17752_o = n17749_o ? 1'b1 : n17751_o;
  /* fpu.vhdl:401:18  */
  assign n17755_o = $unsigned(6'b001110) >= $unsigned(n17663_o);
  assign n17757_o = n17674_o[49];
  /* fpu.vhdl:401:13  */
  assign n17758_o = n17755_o ? 1'b1 : n17757_o;
  /* fpu.vhdl:401:18  */
  assign n17761_o = $unsigned(6'b001111) >= $unsigned(n17663_o);
  assign n17763_o = n17674_o[48];
  /* fpu.vhdl:401:13  */
  assign n17764_o = n17761_o ? 1'b1 : n17763_o;
  /* fpu.vhdl:401:18  */
  assign n17767_o = $unsigned(6'b010000) >= $unsigned(n17663_o);
  assign n17769_o = n17674_o[47];
  /* fpu.vhdl:401:13  */
  assign n17770_o = n17767_o ? 1'b1 : n17769_o;
  /* fpu.vhdl:401:18  */
  assign n17773_o = $unsigned(6'b010001) >= $unsigned(n17663_o);
  assign n17775_o = n17674_o[46];
  /* fpu.vhdl:401:13  */
  assign n17776_o = n17773_o ? 1'b1 : n17775_o;
  /* fpu.vhdl:401:18  */
  assign n17779_o = $unsigned(6'b010010) >= $unsigned(n17663_o);
  assign n17781_o = n17674_o[45];
  /* fpu.vhdl:401:13  */
  assign n17782_o = n17779_o ? 1'b1 : n17781_o;
  /* fpu.vhdl:401:18  */
  assign n17785_o = $unsigned(6'b010011) >= $unsigned(n17663_o);
  assign n17787_o = n17674_o[44];
  /* fpu.vhdl:401:13  */
  assign n17788_o = n17785_o ? 1'b1 : n17787_o;
  /* fpu.vhdl:401:18  */
  assign n17791_o = $unsigned(6'b010100) >= $unsigned(n17663_o);
  assign n17793_o = n17674_o[43];
  /* fpu.vhdl:401:13  */
  assign n17794_o = n17791_o ? 1'b1 : n17793_o;
  /* fpu.vhdl:401:18  */
  assign n17797_o = $unsigned(6'b010101) >= $unsigned(n17663_o);
  assign n17799_o = n17674_o[42];
  /* fpu.vhdl:401:13  */
  assign n17800_o = n17797_o ? 1'b1 : n17799_o;
  /* fpu.vhdl:401:18  */
  assign n17803_o = $unsigned(6'b010110) >= $unsigned(n17663_o);
  assign n17805_o = n17674_o[41];
  /* fpu.vhdl:401:13  */
  assign n17806_o = n17803_o ? 1'b1 : n17805_o;
  /* fpu.vhdl:401:18  */
  assign n17809_o = $unsigned(6'b010111) >= $unsigned(n17663_o);
  assign n17811_o = n17674_o[40];
  /* fpu.vhdl:401:13  */
  assign n17812_o = n17809_o ? 1'b1 : n17811_o;
  /* fpu.vhdl:401:18  */
  assign n17815_o = $unsigned(6'b011000) >= $unsigned(n17663_o);
  assign n17817_o = n17674_o[39];
  /* fpu.vhdl:401:13  */
  assign n17818_o = n17815_o ? 1'b1 : n17817_o;
  /* fpu.vhdl:401:18  */
  assign n17821_o = $unsigned(6'b011001) >= $unsigned(n17663_o);
  assign n17823_o = n17674_o[38];
  /* fpu.vhdl:401:13  */
  assign n17824_o = n17821_o ? 1'b1 : n17823_o;
  /* fpu.vhdl:401:18  */
  assign n17827_o = $unsigned(6'b011010) >= $unsigned(n17663_o);
  assign n17829_o = n17674_o[37];
  /* fpu.vhdl:401:13  */
  assign n17830_o = n17827_o ? 1'b1 : n17829_o;
  /* fpu.vhdl:401:18  */
  assign n17833_o = $unsigned(6'b011011) >= $unsigned(n17663_o);
  assign n17835_o = n17674_o[36];
  /* fpu.vhdl:401:13  */
  assign n17836_o = n17833_o ? 1'b1 : n17835_o;
  /* fpu.vhdl:401:18  */
  assign n17839_o = $unsigned(6'b011100) >= $unsigned(n17663_o);
  assign n17841_o = n17674_o[35];
  /* fpu.vhdl:401:13  */
  assign n17842_o = n17839_o ? 1'b1 : n17841_o;
  /* fpu.vhdl:401:18  */
  assign n17845_o = $unsigned(6'b011101) >= $unsigned(n17663_o);
  assign n17847_o = n17674_o[34];
  /* fpu.vhdl:401:13  */
  assign n17848_o = n17845_o ? 1'b1 : n17847_o;
  /* fpu.vhdl:401:18  */
  assign n17851_o = $unsigned(6'b011110) >= $unsigned(n17663_o);
  assign n17853_o = n17674_o[33];
  /* fpu.vhdl:401:13  */
  assign n17854_o = n17851_o ? 1'b1 : n17853_o;
  /* fpu.vhdl:401:18  */
  assign n17857_o = $unsigned(6'b011111) >= $unsigned(n17663_o);
  assign n17859_o = n17674_o[32];
  /* fpu.vhdl:401:13  */
  assign n17860_o = n17857_o ? 1'b1 : n17859_o;
  /* fpu.vhdl:401:18  */
  assign n17863_o = $unsigned(6'b100000) >= $unsigned(n17663_o);
  assign n17865_o = n17674_o[31];
  /* fpu.vhdl:401:13  */
  assign n17866_o = n17863_o ? 1'b1 : n17865_o;
  /* fpu.vhdl:401:18  */
  assign n17869_o = $unsigned(6'b100001) >= $unsigned(n17663_o);
  assign n17871_o = n17674_o[30];
  /* fpu.vhdl:401:13  */
  assign n17872_o = n17869_o ? 1'b1 : n17871_o;
  /* fpu.vhdl:401:18  */
  assign n17875_o = $unsigned(6'b100010) >= $unsigned(n17663_o);
  assign n17877_o = n17674_o[29];
  /* fpu.vhdl:401:13  */
  assign n17878_o = n17875_o ? 1'b1 : n17877_o;
  /* fpu.vhdl:401:18  */
  assign n17881_o = $unsigned(6'b100011) >= $unsigned(n17663_o);
  assign n17883_o = n17674_o[28];
  /* fpu.vhdl:401:13  */
  assign n17884_o = n17881_o ? 1'b1 : n17883_o;
  /* fpu.vhdl:401:18  */
  assign n17887_o = $unsigned(6'b100100) >= $unsigned(n17663_o);
  assign n17889_o = n17674_o[27];
  /* fpu.vhdl:401:13  */
  assign n17890_o = n17887_o ? 1'b1 : n17889_o;
  /* fpu.vhdl:401:18  */
  assign n17893_o = $unsigned(6'b100101) >= $unsigned(n17663_o);
  assign n17895_o = n17674_o[26];
  /* fpu.vhdl:401:13  */
  assign n17896_o = n17893_o ? 1'b1 : n17895_o;
  /* fpu.vhdl:401:18  */
  assign n17899_o = $unsigned(6'b100110) >= $unsigned(n17663_o);
  assign n17901_o = n17674_o[25];
  /* fpu.vhdl:401:13  */
  assign n17902_o = n17899_o ? 1'b1 : n17901_o;
  /* fpu.vhdl:401:18  */
  assign n17905_o = $unsigned(6'b100111) >= $unsigned(n17663_o);
  assign n17907_o = n17674_o[24];
  /* fpu.vhdl:401:13  */
  assign n17908_o = n17905_o ? 1'b1 : n17907_o;
  /* fpu.vhdl:401:18  */
  assign n17911_o = $unsigned(6'b101000) >= $unsigned(n17663_o);
  assign n17913_o = n17674_o[23];
  /* fpu.vhdl:401:13  */
  assign n17914_o = n17911_o ? 1'b1 : n17913_o;
  /* fpu.vhdl:401:18  */
  assign n17917_o = $unsigned(6'b101001) >= $unsigned(n17663_o);
  assign n17919_o = n17674_o[22];
  /* fpu.vhdl:401:13  */
  assign n17920_o = n17917_o ? 1'b1 : n17919_o;
  /* fpu.vhdl:401:18  */
  assign n17923_o = $unsigned(6'b101010) >= $unsigned(n17663_o);
  assign n17925_o = n17674_o[21];
  /* fpu.vhdl:401:13  */
  assign n17926_o = n17923_o ? 1'b1 : n17925_o;
  /* fpu.vhdl:401:18  */
  assign n17929_o = $unsigned(6'b101011) >= $unsigned(n17663_o);
  assign n17931_o = n17674_o[20];
  /* fpu.vhdl:401:13  */
  assign n17932_o = n17929_o ? 1'b1 : n17931_o;
  /* fpu.vhdl:401:18  */
  assign n17935_o = $unsigned(6'b101100) >= $unsigned(n17663_o);
  assign n17937_o = n17674_o[19];
  /* fpu.vhdl:401:13  */
  assign n17938_o = n17935_o ? 1'b1 : n17937_o;
  /* fpu.vhdl:401:18  */
  assign n17941_o = $unsigned(6'b101101) >= $unsigned(n17663_o);
  assign n17943_o = n17674_o[18];
  /* fpu.vhdl:401:13  */
  assign n17944_o = n17941_o ? 1'b1 : n17943_o;
  /* fpu.vhdl:401:18  */
  assign n17947_o = $unsigned(6'b101110) >= $unsigned(n17663_o);
  assign n17949_o = n17674_o[17];
  /* fpu.vhdl:401:13  */
  assign n17950_o = n17947_o ? 1'b1 : n17949_o;
  /* fpu.vhdl:401:18  */
  assign n17953_o = $unsigned(6'b101111) >= $unsigned(n17663_o);
  assign n17955_o = n17674_o[16];
  /* fpu.vhdl:401:13  */
  assign n17956_o = n17953_o ? 1'b1 : n17955_o;
  /* fpu.vhdl:401:18  */
  assign n17959_o = $unsigned(6'b110000) >= $unsigned(n17663_o);
  assign n17961_o = n17674_o[15];
  /* fpu.vhdl:401:13  */
  assign n17962_o = n17959_o ? 1'b1 : n17961_o;
  /* fpu.vhdl:401:18  */
  assign n17965_o = $unsigned(6'b110001) >= $unsigned(n17663_o);
  assign n17967_o = n17674_o[14];
  /* fpu.vhdl:401:13  */
  assign n17968_o = n17965_o ? 1'b1 : n17967_o;
  /* fpu.vhdl:401:18  */
  assign n17971_o = $unsigned(6'b110010) >= $unsigned(n17663_o);
  assign n17973_o = n17674_o[13];
  /* fpu.vhdl:401:13  */
  assign n17974_o = n17971_o ? 1'b1 : n17973_o;
  /* fpu.vhdl:401:18  */
  assign n17977_o = $unsigned(6'b110011) >= $unsigned(n17663_o);
  assign n17979_o = n17674_o[12];
  /* fpu.vhdl:401:13  */
  assign n17980_o = n17977_o ? 1'b1 : n17979_o;
  /* fpu.vhdl:401:18  */
  assign n17983_o = $unsigned(6'b110100) >= $unsigned(n17663_o);
  assign n17985_o = n17674_o[11];
  /* fpu.vhdl:401:13  */
  assign n17986_o = n17983_o ? 1'b1 : n17985_o;
  /* fpu.vhdl:401:18  */
  assign n17989_o = $unsigned(6'b110101) >= $unsigned(n17663_o);
  assign n17991_o = n17674_o[10];
  /* fpu.vhdl:401:13  */
  assign n17992_o = n17989_o ? 1'b1 : n17991_o;
  /* fpu.vhdl:401:18  */
  assign n17995_o = $unsigned(6'b110110) >= $unsigned(n17663_o);
  assign n17997_o = n17674_o[9];
  /* fpu.vhdl:401:13  */
  assign n17998_o = n17995_o ? 1'b1 : n17997_o;
  /* fpu.vhdl:401:18  */
  assign n18001_o = $unsigned(6'b110111) >= $unsigned(n17663_o);
  assign n18003_o = n17674_o[8];
  /* fpu.vhdl:401:13  */
  assign n18004_o = n18001_o ? 1'b1 : n18003_o;
  /* fpu.vhdl:401:18  */
  assign n18007_o = $unsigned(6'b111000) >= $unsigned(n17663_o);
  assign n18009_o = n17674_o[7];
  /* fpu.vhdl:401:13  */
  assign n18010_o = n18007_o ? 1'b1 : n18009_o;
  /* fpu.vhdl:401:18  */
  assign n18013_o = $unsigned(6'b111001) >= $unsigned(n17663_o);
  assign n18015_o = n17674_o[6];
  /* fpu.vhdl:401:13  */
  assign n18016_o = n18013_o ? 1'b1 : n18015_o;
  /* fpu.vhdl:401:18  */
  assign n18019_o = $unsigned(6'b111010) >= $unsigned(n17663_o);
  assign n18021_o = n17674_o[5];
  /* fpu.vhdl:401:13  */
  assign n18022_o = n18019_o ? 1'b1 : n18021_o;
  /* fpu.vhdl:401:18  */
  assign n18025_o = $unsigned(6'b111011) >= $unsigned(n17663_o);
  assign n18027_o = n17674_o[4];
  /* fpu.vhdl:401:13  */
  assign n18028_o = n18025_o ? 1'b1 : n18027_o;
  /* fpu.vhdl:401:18  */
  assign n18031_o = $unsigned(6'b111100) >= $unsigned(n17663_o);
  assign n18033_o = n17674_o[3];
  /* fpu.vhdl:401:13  */
  assign n18034_o = n18031_o ? 1'b1 : n18033_o;
  /* fpu.vhdl:401:18  */
  assign n18037_o = $unsigned(6'b111101) >= $unsigned(n17663_o);
  assign n18039_o = n17674_o[2];
  /* fpu.vhdl:401:13  */
  assign n18040_o = n18037_o ? 1'b1 : n18039_o;
  /* fpu.vhdl:401:18  */
  assign n18043_o = $unsigned(6'b111110) >= $unsigned(n17663_o);
  assign n18045_o = n17674_o[1];
  /* fpu.vhdl:401:13  */
  assign n18046_o = n18043_o ? 1'b1 : n18045_o;
  assign n18047_o = n17674_o[0];
  /* fpu.vhdl:401:18  */
  assign n18049_o = $unsigned(6'b111111) >= $unsigned(n17663_o);
  /* fpu.vhdl:401:13  */
  assign n18051_o = n18049_o ? 1'b1 : n18047_o;
  assign n18052_o = {n17673_o, n17680_o, n17686_o, n17692_o, n17698_o, n17704_o, n17710_o, n17716_o, n17722_o, n17728_o, n17734_o, n17740_o, n17746_o, n17752_o, n17758_o, n17764_o, n17770_o, n17776_o, n17782_o, n17788_o, n17794_o, n17800_o, n17806_o, n17812_o, n17818_o, n17824_o, n17830_o, n17836_o, n17842_o, n17848_o, n17854_o, n17860_o, n17866_o, n17872_o, n17878_o, n17884_o, n17890_o, n17896_o, n17902_o, n17908_o, n17914_o, n17920_o, n17926_o, n17932_o, n17938_o, n17944_o, n17950_o, n17956_o, n17962_o, n17968_o, n17974_o, n17980_o, n17986_o, n17992_o, n17998_o, n18004_o, n18010_o, n18016_o, n18022_o, n18028_o, n18034_o, n18040_o, n18046_o, n18051_o};
  /* fpu.vhdl:2378:9  */
  assign n18054_o = n17661_o ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n18052_o;
  /* fpu.vhdl:2376:9  */
  assign n18056_o = n17659_o ? 64'b1111111111111111111111111111111111111111111111111111111111111111 : n18054_o;
  /* fpu.vhdl:2383:16  */
  assign n18057_o = r[715:714];
  /* fpu.vhdl:2385:28  */
  assign n18058_o = r[462:399];
  /* fpu.vhdl:2384:13  */
  assign n18060_o = n18057_o == 2'b00;
  /* fpu.vhdl:2387:28  */
  assign n18061_o = r[238:159];
  /* fpu.vhdl:2387:30  */
  assign n18062_o = n18061_o[79:16];
  /* fpu.vhdl:2386:13  */
  assign n18064_o = n18057_o == 2'b01;
  /* fpu.vhdl:2389:28  */
  assign n18065_o = r[318:239];
  /* fpu.vhdl:2389:30  */
  assign n18066_o = n18065_o[79:16];
  /* fpu.vhdl:2388:13  */
  assign n18068_o = n18057_o == 2'b10;
  /* fpu.vhdl:2391:28  */
  assign n18069_o = r[398:319];
  /* fpu.vhdl:2391:30  */
  assign n18070_o = n18069_o[79:16];
  assign n18071_o = {n18068_o, n18064_o, n18060_o};
  /* fpu.vhdl:2383:9  */
  always @*
    case (n18071_o)
      3'b100: n18072_o = n18066_o;
      3'b010: n18072_o = n18062_o;
      3'b001: n18072_o = n18058_o;
      default: n18072_o = n18070_o;
    endcase
  /* fpu.vhdl:2393:22  */
  assign n18073_o = n18056_o & n18072_o;
  /* fpu.vhdl:2393:13  */
  assign n18074_o = |(n18073_o);
  /* fpu.vhdl:2393:40  */
  assign n18075_o = n18074_o & n17442_o;
  /* fpu.vhdl:2393:9  */
  assign n18077_o = n18075_o ? 1'b1 : n17157_o;
  /* fpu.vhdl:2397:22  */
  assign n18078_o = ~n18072_o;
  /* fpu.vhdl:2396:9  */
  assign n18079_o = opsel_ainv ? n18078_o : n18072_o;
  /* fpu.vhdl:2401:13  */
  assign n18081_o = opsel_b == 2'b00;
  /* fpu.vhdl:2404:28  */
  assign n18082_o = r[462:399];
  /* fpu.vhdl:2403:13  */
  assign n18084_o = opsel_b == 2'b01;
  /* fpu.vhdl:2406:39  */
  assign n18085_o = r[126];
  /* fpu.vhdl:2406:63  */
  assign n18086_o = r[126];
  /* fpu.vhdl:2406:57  */
  assign n18087_o = ~n18086_o;
  assign n18150_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18151_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18152_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18153_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18154_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18155_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18156_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18157_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18158_o = {n18085_o, 1'b0, 1'b0, 1'b0};
  assign n18159_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18160_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18161_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18162_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18163_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18164_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n18165_o = {1'b0, n18087_o, 1'b0, 1'b0};
  assign n18166_o = {n18150_o, n18151_o, n18152_o, n18153_o};
  assign n18167_o = {n18154_o, n18155_o, n18156_o, n18157_o};
  assign n18168_o = {n18158_o, n18159_o, n18160_o, n18161_o};
  assign n18169_o = {n18162_o, n18163_o, n18164_o, n18165_o};
  assign n18170_o = {n18166_o, n18167_o, n18168_o, n18169_o};
  /* fpu.vhdl:2405:13  */
  assign n18172_o = opsel_b == 2'b10;
  /* fpu.vhdl:2410:61  */
  assign n18173_o = r[527:522];
  /* fpu.vhdl:2410:44  */
  assign n18174_o = {{58{n18173_o[5]}}, n18173_o}; // sext
  assign n18175_o = {n18172_o, n18084_o, n18081_o};
  /* fpu.vhdl:2400:9  */
  always @*
    case (n18175_o)
      3'b100: n18177_o = n18170_o;
      3'b010: n18177_o = n18082_o;
      3'b001: n18177_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      default: n18177_o = n18174_o;
    endcase
  /* fpu.vhdl:2413:22  */
  assign n18179_o = ~n18177_o;
  /* fpu.vhdl:2412:9  */
  assign n18180_o = opsel_binv ? n18179_o : n18177_o;
  /* fpu.vhdl:2416:14  */
  assign n18181_o = r[676:664];
  /* fpu.vhdl:2416:20  */
  assign n18183_o = $signed(n18181_o) >= $signed(13'b1111111000000);
  /* fpu.vhdl:2416:54  */
  assign n18184_o = r[676:664];
  /* fpu.vhdl:2416:60  */
  assign n18186_o = $signed(n18184_o) <= $signed(13'b0000000111111);
  /* fpu.vhdl:2416:48  */
  assign n18187_o = n18183_o & n18186_o;
  /* fpu.vhdl:2417:39  */
  assign n18189_o = r[462:399];
  /* fpu.vhdl:2417:58  */
  assign n18190_o = r[518];
  /* fpu.vhdl:2417:52  */
  assign n18191_o = n17504_o | n18190_o;
  /* fpu.vhdl:2417:41  */
  assign n18192_o = {n18189_o, n18191_o};
  /* fpu.vhdl:2417:69  */
  assign n18193_o = r[517:463];
  /* fpu.vhdl:2417:64  */
  assign n18194_o = {n18192_o, n18193_o};
  /* fpu.vhdl:2418:62  */
  assign n18195_o = r[670:664];
  /* fpu.vhdl:351:19  */
  assign n18203_o = n18195_o[6:5];
  /* fpu.vhdl:353:26  */
  assign n18204_o = n18194_o[119:25];
  /* fpu.vhdl:352:13  */
  assign n18206_o = n18203_o == 2'b00;
  /* fpu.vhdl:355:26  */
  assign n18207_o = n18194_o[87:0];
  /* fpu.vhdl:355:40  */
  assign n18209_o = {n18207_o, 7'b0000000};
  /* fpu.vhdl:354:13  */
  assign n18211_o = n18203_o == 2'b01;
  /* fpu.vhdl:357:48  */
  assign n18212_o = n18194_o[119:89];
  /* fpu.vhdl:357:43  */
  assign n18214_o = {64'b0000000000000000000000000000000000000000000000000000000000000000, n18212_o};
  /* fpu.vhdl:356:13  */
  assign n18216_o = n18203_o == 2'b10;
  /* fpu.vhdl:359:40  */
  assign n18217_o = n18194_o[119:57];
  /* fpu.vhdl:359:35  */
  assign n18219_o = {32'b00000000000000000000000000000000, n18217_o};
  assign n18220_o = {n18216_o, n18211_o, n18206_o};
  /* fpu.vhdl:351:9  */
  always @*
    case (n18220_o)
      3'b100: n18221_o = n18214_o;
      3'b010: n18221_o = n18209_o;
      3'b001: n18221_o = n18204_o;
      default: n18221_o = n18219_o;
    endcase
  /* fpu.vhdl:361:19  */
  assign n18223_o = n18195_o[4:3];
  /* fpu.vhdl:363:25  */
  assign n18224_o = n18221_o[94:24];
  /* fpu.vhdl:362:13  */
  assign n18226_o = n18223_o == 2'b00;
  /* fpu.vhdl:365:25  */
  assign n18227_o = n18221_o[86:16];
  /* fpu.vhdl:364:13  */
  assign n18229_o = n18223_o == 2'b01;
  /* fpu.vhdl:367:25  */
  assign n18230_o = n18221_o[78:8];
  /* fpu.vhdl:366:13  */
  assign n18232_o = n18223_o == 2'b10;
  /* fpu.vhdl:369:25  */
  assign n18233_o = n18221_o[70:0];
  assign n18234_o = {n18232_o, n18229_o, n18226_o};
  /* fpu.vhdl:361:9  */
  always @*
    case (n18234_o)
      3'b100: n18235_o = n18230_o;
      3'b010: n18235_o = n18227_o;
      3'b001: n18235_o = n18224_o;
      default: n18235_o = n18233_o;
    endcase
  /* fpu.vhdl:371:19  */
  assign n18237_o = n18195_o[2:0];
  /* fpu.vhdl:373:29  */
  assign n18238_o = n18235_o[70:7];
  /* fpu.vhdl:372:13  */
  assign n18240_o = n18237_o == 3'b000;
  /* fpu.vhdl:375:29  */
  assign n18241_o = n18235_o[69:6];
  /* fpu.vhdl:374:13  */
  assign n18243_o = n18237_o == 3'b001;
  /* fpu.vhdl:377:29  */
  assign n18244_o = n18235_o[68:5];
  /* fpu.vhdl:376:13  */
  assign n18246_o = n18237_o == 3'b010;
  /* fpu.vhdl:379:29  */
  assign n18247_o = n18235_o[67:4];
  /* fpu.vhdl:378:13  */
  assign n18249_o = n18237_o == 3'b011;
  /* fpu.vhdl:381:29  */
  assign n18250_o = n18235_o[66:3];
  /* fpu.vhdl:380:13  */
  assign n18252_o = n18237_o == 3'b100;
  /* fpu.vhdl:383:29  */
  assign n18253_o = n18235_o[65:2];
  /* fpu.vhdl:382:13  */
  assign n18255_o = n18237_o == 3'b101;
  /* fpu.vhdl:385:29  */
  assign n18256_o = n18235_o[64:1];
  /* fpu.vhdl:384:13  */
  assign n18258_o = n18237_o == 3'b110;
  /* fpu.vhdl:387:29  */
  assign n18259_o = n18235_o[63:0];
  assign n18260_o = {n18258_o, n18255_o, n18252_o, n18249_o, n18246_o, n18243_o, n18240_o};
  /* fpu.vhdl:371:9  */
  always @*
    case (n18260_o)
      7'b1000000: n18261_o = n18256_o;
      7'b0100000: n18261_o = n18253_o;
      7'b0010000: n18261_o = n18250_o;
      7'b0001000: n18261_o = n18247_o;
      7'b0000100: n18261_o = n18244_o;
      7'b0000010: n18261_o = n18241_o;
      7'b0000001: n18261_o = n18238_o;
      default: n18261_o = n18259_o;
    endcase
  /* fpu.vhdl:2416:9  */
  assign n18264_o = n18187_o ? n18261_o : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* fpu.vhdl:2422:49  */
  assign n18265_o = in_a + in_b;
  /* fpu.vhdl:2422:66  */
  assign n18266_o = {63'b0, carry_in};  //  uext
  /* fpu.vhdl:2422:66  */
  assign n18267_o = n18265_o + n18266_o;
  /* fpu.vhdl:2425:18  */
  assign n18269_o = r[126];
  assign n18271_o = n18267_o[30:2];
  /* fpu.vhdl:2425:13  */
  assign n18272_o = n18269_o ? 29'b00000000000000000000000000000 : n18271_o;
  assign n18273_o = {n18272_o, 2'b00};
  assign n18274_o = n18267_o[30:0];
  /* fpu.vhdl:2423:9  */
  assign n18275_o = opsel_mask ? n18273_o : n18274_o;
  assign n18276_o = n18267_o[63:31];
  assign n18277_o = {n18276_o, n18275_o};
  /* fpu.vhdl:2430:13  */
  assign n18279_o = opsel_r == 2'b00;
  /* fpu.vhdl:2432:13  */
  assign n18281_o = opsel_r == 2'b01;
  /* fpu.vhdl:2435:47  */
  assign n18282_o = multiply_to_f[122:59];
  /* fpu.vhdl:2434:13  */
  assign n18284_o = opsel_r == 2'b10;
  /* fpu.vhdl:2439:50  */
  assign n18285_o = r[158:127];
  assign n18286_o = {n17382_o, n17378_o, n17374_o, n17370_o, n17366_o, n17362_o, n17358_o, n17354_o};
  /* fpu.vhdl:2439:56  */
  assign n18287_o = n18285_o & n18286_o;
  /* fpu.vhdl:2439:45  */
  assign n18289_o = {32'b00000000000000000000000000000000, n18287_o};
  /* fpu.vhdl:2438:21  */
  assign n18291_o = misc_sel == 4'b0000;
  /* fpu.vhdl:2440:21  */
  assign n18293_o = misc_sel == 4'b0001;
  /* fpu.vhdl:2443:21  */
  assign n18295_o = misc_sel == 4'b0010;
  /* fpu.vhdl:2446:21  */
  assign n18297_o = misc_sel == 4'b0011;
  /* fpu.vhdl:2451:45  */
  assign n18298_o = r[206:175];
  /* fpu.vhdl:2451:73  */
  assign n18299_o = r[286:255];
  /* fpu.vhdl:2451:59  */
  assign n18300_o = {n18298_o, n18299_o};
  /* fpu.vhdl:2449:21  */
  assign n18302_o = misc_sel == 4'b0100;
  /* fpu.vhdl:2454:45  */
  assign n18303_o = r[238:207];
  /* fpu.vhdl:2454:74  */
  assign n18304_o = r[318:287];
  /* fpu.vhdl:2454:60  */
  assign n18305_o = {n18303_o, n18304_o};
  /* fpu.vhdl:2452:21  */
  assign n18307_o = misc_sel == 4'b0110;
  /* fpu.vhdl:2456:42  */
  assign n18309_o = {10'b0000000000, inverse_est};
  /* fpu.vhdl:2456:56  */
  assign n18311_o = {n18309_o, 35'b00000000000000000000000000000000000};
  /* fpu.vhdl:2455:21  */
  assign n18313_o = misc_sel == 4'b0111;
  /* fpu.vhdl:2457:21  */
  assign n18315_o = misc_sel == 4'b1000;
  /* fpu.vhdl:2460:21  */
  assign n18317_o = misc_sel == 4'b1001;
  /* fpu.vhdl:2463:21  */
  assign n18319_o = misc_sel == 4'b1010;
  /* fpu.vhdl:2466:21  */
  assign n18321_o = misc_sel == 4'b1011;
  /* fpu.vhdl:2469:21  */
  assign n18323_o = misc_sel == 4'b1100;
  /* fpu.vhdl:2472:21  */
  assign n18325_o = misc_sel == 4'b1101;
  /* fpu.vhdl:2475:21  */
  assign n18327_o = misc_sel == 4'b1110;
  /* fpu.vhdl:2478:21  */
  assign n18329_o = misc_sel == 4'b1111;
  assign n18330_o = {n18329_o, n18327_o, n18325_o, n18323_o, n18321_o, n18319_o, n18317_o, n18315_o, n18313_o, n18307_o, n18302_o, n18297_o, n18295_o, n18293_o, n18291_o};
  /* fpu.vhdl:2437:17  */
  always @*
    case (n18330_o)
      15'b100000000000000: n18343_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      15'b010000000000000: n18343_o = 64'b1111111111111111111111111111111111111111111111111111111111111111;
      15'b001000000000000: n18343_o = 64'b1000000000000000000000000000000000000000000000000000000000000000;
      15'b000100000000000: n18343_o = 64'b0111111111111111111111111111111111111111111111111111111111111111;
      15'b000010000000000: n18343_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      15'b000001000000000: n18343_o = 64'b0000000000000000000000000000000011111111111111111111111111111111;
      15'b000000100000000: n18343_o = 64'b1111111111111111111111111111111110000000000000000000000000000000;
      15'b000000010000000: n18343_o = 64'b0000000000000000000000000000000001111111111111111111111111111111;
      15'b000000001000000: n18343_o = n18311_o;
      15'b000000000100000: n18343_o = n18305_o;
      15'b000000000010000: n18343_o = n18300_o;
      15'b000000000001000: n18343_o = 64'b0000000001111111111111111111111110000000000000000000000000000000;
      15'b000000000000100: n18343_o = 64'b0000000001111111111111111111111111111111111111111111111111111100;
      15'b000000000000010: n18343_o = 64'b0000000000100000000000000000000000000000000000000000000000000000;
      15'b000000000000001: n18343_o = n18289_o;
      default: n18343_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    endcase
  assign n18344_o = {n18284_o, n18281_o, n18279_o};
  /* fpu.vhdl:2429:9  */
  always @*
    case (n18344_o)
      3'b100: n18345_o = n18282_o;
      3'b010: n18345_o = n18264_o;
      3'b001: n18345_o = n18277_o;
      default: n18345_o = n18343_o;
    endcase
  assign n18347_o = r[518:463];
  /* fpu.vhdl:2490:61  */
  assign n18348_o = r[518:463];
  /* fpu.vhdl:2490:55  */
  assign n18349_o = ~n18348_o;
  /* fpu.vhdl:2490:73  */
  assign n18350_o = r[519];
  /* fpu.vhdl:2490:67  */
  assign n18351_o = ~n18350_o;
  /* fpu.vhdl:2490:64  */
  assign n18352_o = {55'b0, n18351_o};  //  uext
  /* fpu.vhdl:2490:64  */
  assign n18353_o = n18349_o + n18352_o;
  /* fpu.vhdl:2489:17  */
  assign n18355_o = opsel_s == 2'b01;
  /* fpu.vhdl:2492:48  */
  assign n18356_o = multiply_to_f[58:3];
  /* fpu.vhdl:2491:17  */
  assign n18358_o = opsel_s == 2'b11;
  /* fpu.vhdl:2494:37  */
  assign n18359_o = n18264_o[63:8];
  /* fpu.vhdl:2495:33  */
  assign n18360_o = n18264_o[7:0];
  /* fpu.vhdl:2495:46  */
  assign n18362_o = n18360_o != 8'b00000000;
  /* fpu.vhdl:2495:21  */
  assign n18364_o = n18362_o ? 1'b1 : n18077_o;
  /* fpu.vhdl:2493:17  */
  assign n18366_o = opsel_s == 2'b10;
  assign n18368_o = {n18366_o, n18358_o, n18355_o};
  /* fpu.vhdl:2488:13  */
  always @*
    case (n18368_o)
      3'b100: n18369_o = n18359_o;
      3'b010: n18369_o = n18356_o;
      3'b001: n18369_o = n18353_o;
      default: n18369_o = 56'b00000000000000000000000000000000000000000000000000000000;
    endcase
  /* fpu.vhdl:2488:13  */
  always @*
    case (n18368_o)
      3'b100: n18370_o = n18364_o;
      3'b010: n18370_o = n18077_o;
      3'b001: n18370_o = n18077_o;
      default: n18370_o = n18077_o;
    endcase
  assign n18371_o = {n18370_o, n18369_o};
  assign n18372_o = {n18077_o, n18347_o};
  /* fpu.vhdl:2487:9  */
  assign n18373_o = n17476_o ? n18371_o : n18372_o;
  assign n18374_o = {n18264_o, n13526_o};
  assign n18375_o = n13464_o[79:3];
  assign n18376_o = r[238:162];
  /* fpu.vhdl:650:9  */
  assign n18377_o = n13152_o ? n18375_o : n18376_o;
  /* fpu.vhdl:2503:9  */
  assign n18378_o = n17454_o ? n18374_o : n18377_o;
  assign n18382_o = n13464_o[2:0];
  assign n18383_o = r[161:159];
  /* fpu.vhdl:650:9  */
  assign n18384_o = n13152_o ? n18382_o : n18383_o;
  assign n18385_o = {n18264_o, n13526_o};
  assign n18386_o = n13464_o[159:83];
  assign n18387_o = r[318:242];
  /* fpu.vhdl:650:9  */
  assign n18388_o = n13152_o ? n18386_o : n18387_o;
  /* fpu.vhdl:2507:9  */
  assign n18389_o = n17459_o ? n18385_o : n18388_o;
  assign n18393_o = n13464_o[82:80];
  assign n18394_o = r[241:239];
  /* fpu.vhdl:650:9  */
  assign n18395_o = n13152_o ? n18393_o : n18394_o;
  assign n18396_o = {n18264_o, n13526_o};
  assign n18397_o = n13464_o[239:163];
  assign n18398_o = r[398:322];
  /* fpu.vhdl:650:9  */
  assign n18399_o = n13152_o ? n18397_o : n18398_o;
  /* fpu.vhdl:2511:9  */
  assign n18400_o = n17464_o ? n18396_o : n18399_o;
  assign n18401_o = n13464_o[162:160];
  assign n18402_o = r[321:319];
  /* fpu.vhdl:650:9  */
  assign n18403_o = n13152_o ? n18401_o : n18402_o;
  /* fpu.vhdl:2516:20  */
  assign n18405_o = opsel_r == 2'b01;
  /* fpu.vhdl:2516:9  */
  assign n18406_o = n18405_o ? n13526_o : n17171_o;
  /* fpu.vhdl:2521:40  */
  assign n18408_o = r[462:399];
  /* helpers.vhdl:221:43  */
  assign n18420_o = n18408_o[0];
  /* helpers.vhdl:221:43  */
  assign n18423_o = n18408_o[1];
  /* helpers.vhdl:221:43  */
  assign n18425_o = n18408_o[2];
  /* helpers.vhdl:221:43  */
  assign n18427_o = n18408_o[3];
  /* helpers.vhdl:221:43  */
  assign n18429_o = n18408_o[4];
  /* helpers.vhdl:221:43  */
  assign n18431_o = n18408_o[5];
  /* helpers.vhdl:221:43  */
  assign n18433_o = n18408_o[6];
  /* helpers.vhdl:221:43  */
  assign n18435_o = n18408_o[7];
  /* helpers.vhdl:221:43  */
  assign n18437_o = n18408_o[8];
  /* helpers.vhdl:221:43  */
  assign n18439_o = n18408_o[9];
  /* helpers.vhdl:221:43  */
  assign n18441_o = n18408_o[10];
  /* helpers.vhdl:221:43  */
  assign n18443_o = n18408_o[11];
  /* helpers.vhdl:221:43  */
  assign n18445_o = n18408_o[12];
  /* helpers.vhdl:221:43  */
  assign n18447_o = n18408_o[13];
  /* helpers.vhdl:221:43  */
  assign n18449_o = n18408_o[14];
  /* helpers.vhdl:221:43  */
  assign n18451_o = n18408_o[15];
  /* helpers.vhdl:221:43  */
  assign n18453_o = n18408_o[16];
  /* helpers.vhdl:221:43  */
  assign n18455_o = n18408_o[17];
  /* helpers.vhdl:221:43  */
  assign n18457_o = n18408_o[18];
  /* helpers.vhdl:221:43  */
  assign n18459_o = n18408_o[19];
  /* helpers.vhdl:221:43  */
  assign n18461_o = n18408_o[20];
  /* helpers.vhdl:221:43  */
  assign n18463_o = n18408_o[21];
  /* helpers.vhdl:221:43  */
  assign n18465_o = n18408_o[22];
  /* helpers.vhdl:221:43  */
  assign n18467_o = n18408_o[23];
  /* helpers.vhdl:221:43  */
  assign n18469_o = n18408_o[24];
  /* helpers.vhdl:221:43  */
  assign n18471_o = n18408_o[25];
  /* helpers.vhdl:221:43  */
  assign n18473_o = n18408_o[26];
  /* helpers.vhdl:221:43  */
  assign n18475_o = n18408_o[27];
  /* helpers.vhdl:221:43  */
  assign n18477_o = n18408_o[28];
  /* helpers.vhdl:221:43  */
  assign n18479_o = n18408_o[29];
  /* helpers.vhdl:221:43  */
  assign n18481_o = n18408_o[30];
  /* helpers.vhdl:221:43  */
  assign n18483_o = n18408_o[31];
  /* helpers.vhdl:221:43  */
  assign n18485_o = n18408_o[32];
  /* helpers.vhdl:221:43  */
  assign n18487_o = n18408_o[33];
  /* helpers.vhdl:221:43  */
  assign n18489_o = n18408_o[34];
  /* helpers.vhdl:221:43  */
  assign n18491_o = n18408_o[35];
  /* helpers.vhdl:221:43  */
  assign n18493_o = n18408_o[36];
  /* helpers.vhdl:221:43  */
  assign n18495_o = n18408_o[37];
  /* helpers.vhdl:221:43  */
  assign n18497_o = n18408_o[38];
  /* helpers.vhdl:221:43  */
  assign n18499_o = n18408_o[39];
  /* helpers.vhdl:221:43  */
  assign n18501_o = n18408_o[40];
  /* helpers.vhdl:221:43  */
  assign n18503_o = n18408_o[41];
  /* helpers.vhdl:221:43  */
  assign n18505_o = n18408_o[42];
  /* helpers.vhdl:221:43  */
  assign n18507_o = n18408_o[43];
  /* helpers.vhdl:221:43  */
  assign n18509_o = n18408_o[44];
  /* helpers.vhdl:221:43  */
  assign n18511_o = n18408_o[45];
  /* helpers.vhdl:221:43  */
  assign n18513_o = n18408_o[46];
  /* helpers.vhdl:221:43  */
  assign n18515_o = n18408_o[47];
  /* helpers.vhdl:221:43  */
  assign n18517_o = n18408_o[48];
  /* helpers.vhdl:221:43  */
  assign n18519_o = n18408_o[49];
  /* helpers.vhdl:221:43  */
  assign n18521_o = n18408_o[50];
  /* helpers.vhdl:221:43  */
  assign n18523_o = n18408_o[51];
  /* helpers.vhdl:221:43  */
  assign n18525_o = n18408_o[52];
  /* helpers.vhdl:221:43  */
  assign n18527_o = n18408_o[53];
  /* helpers.vhdl:221:43  */
  assign n18529_o = n18408_o[54];
  /* helpers.vhdl:221:43  */
  assign n18531_o = n18408_o[55];
  /* helpers.vhdl:221:43  */
  assign n18533_o = n18408_o[56];
  /* helpers.vhdl:221:43  */
  assign n18535_o = n18408_o[57];
  /* helpers.vhdl:221:43  */
  assign n18537_o = n18408_o[58];
  /* helpers.vhdl:221:43  */
  assign n18539_o = n18408_o[59];
  /* helpers.vhdl:221:43  */
  assign n18541_o = n18408_o[60];
  /* helpers.vhdl:221:43  */
  assign n18543_o = n18408_o[61];
  /* helpers.vhdl:221:43  */
  assign n18545_o = n18408_o[62];
  /* helpers.vhdl:221:43  */
  assign n18547_o = n18408_o[63];
  assign n18548_o = {n18420_o, n18423_o, n18425_o, n18427_o, n18429_o, n18431_o, n18433_o, n18435_o, n18437_o, n18439_o, n18441_o, n18443_o, n18445_o, n18447_o, n18449_o, n18451_o, n18453_o, n18455_o, n18457_o, n18459_o, n18461_o, n18463_o, n18465_o, n18467_o, n18469_o, n18471_o, n18473_o, n18475_o, n18477_o, n18479_o, n18481_o, n18483_o, n18485_o, n18487_o, n18489_o, n18491_o, n18493_o, n18495_o, n18497_o, n18499_o, n18501_o, n18503_o, n18505_o, n18507_o, n18509_o, n18511_o, n18513_o, n18515_o, n18517_o, n18519_o, n18521_o, n18523_o, n18525_o, n18527_o, n18529_o, n18531_o, n18533_o, n18535_o, n18537_o, n18539_o, n18541_o, n18543_o, n18545_o, n18547_o};
  /* helpers.vhdl:282:34  */
  assign n18561_o = -n18548_o;
  /* helpers.vhdl:283:23  */
  assign n18563_o = n18561_o & n18548_o;
  /* helpers.vhdl:284:21  */
  assign n18565_o = n18561_o | n18548_o;
  /* helpers.vhdl:266:29  */
  assign n18576_o = n18565_o[1];
  /* helpers.vhdl:266:55  */
  assign n18577_o = n18565_o[0];
  /* helpers.vhdl:266:50  */
  assign n18578_o = ~n18577_o;
  /* helpers.vhdl:266:46  */
  assign n18579_o = n18576_o & n18578_o;
  /* helpers.vhdl:266:24  */
  assign n18581_o = 1'b0 | n18579_o;
  /* helpers.vhdl:266:29  */
  assign n18583_o = n18565_o[3];
  /* helpers.vhdl:266:55  */
  assign n18584_o = n18565_o[2];
  /* helpers.vhdl:266:50  */
  assign n18585_o = ~n18584_o;
  /* helpers.vhdl:266:46  */
  assign n18586_o = n18583_o & n18585_o;
  /* helpers.vhdl:266:24  */
  assign n18587_o = n18581_o | n18586_o;
  /* helpers.vhdl:266:29  */
  assign n18588_o = n18565_o[5];
  /* helpers.vhdl:266:55  */
  assign n18589_o = n18565_o[4];
  /* helpers.vhdl:266:50  */
  assign n18590_o = ~n18589_o;
  /* helpers.vhdl:266:46  */
  assign n18591_o = n18588_o & n18590_o;
  /* helpers.vhdl:266:24  */
  assign n18592_o = n18587_o | n18591_o;
  /* helpers.vhdl:266:29  */
  assign n18593_o = n18565_o[7];
  /* helpers.vhdl:266:55  */
  assign n18594_o = n18565_o[6];
  /* helpers.vhdl:266:50  */
  assign n18595_o = ~n18594_o;
  /* helpers.vhdl:266:46  */
  assign n18596_o = n18593_o & n18595_o;
  /* helpers.vhdl:266:24  */
  assign n18597_o = n18592_o | n18596_o;
  /* helpers.vhdl:266:29  */
  assign n18598_o = n18565_o[9];
  /* helpers.vhdl:266:55  */
  assign n18599_o = n18565_o[8];
  /* helpers.vhdl:266:50  */
  assign n18600_o = ~n18599_o;
  /* helpers.vhdl:266:46  */
  assign n18601_o = n18598_o & n18600_o;
  /* helpers.vhdl:266:24  */
  assign n18602_o = n18597_o | n18601_o;
  /* helpers.vhdl:266:29  */
  assign n18603_o = n18565_o[11];
  /* helpers.vhdl:266:55  */
  assign n18604_o = n18565_o[10];
  /* helpers.vhdl:266:50  */
  assign n18605_o = ~n18604_o;
  /* helpers.vhdl:266:46  */
  assign n18606_o = n18603_o & n18605_o;
  /* helpers.vhdl:266:24  */
  assign n18607_o = n18602_o | n18606_o;
  /* helpers.vhdl:266:29  */
  assign n18608_o = n18565_o[13];
  /* helpers.vhdl:266:55  */
  assign n18609_o = n18565_o[12];
  /* helpers.vhdl:266:50  */
  assign n18610_o = ~n18609_o;
  /* helpers.vhdl:266:46  */
  assign n18611_o = n18608_o & n18610_o;
  /* helpers.vhdl:266:24  */
  assign n18612_o = n18607_o | n18611_o;
  /* helpers.vhdl:266:29  */
  assign n18613_o = n18565_o[15];
  /* helpers.vhdl:266:55  */
  assign n18614_o = n18565_o[14];
  /* helpers.vhdl:266:50  */
  assign n18615_o = ~n18614_o;
  /* helpers.vhdl:266:46  */
  assign n18616_o = n18613_o & n18615_o;
  /* helpers.vhdl:266:24  */
  assign n18617_o = n18612_o | n18616_o;
  /* helpers.vhdl:266:29  */
  assign n18618_o = n18565_o[17];
  /* helpers.vhdl:266:55  */
  assign n18619_o = n18565_o[16];
  /* helpers.vhdl:266:50  */
  assign n18620_o = ~n18619_o;
  /* helpers.vhdl:266:46  */
  assign n18621_o = n18618_o & n18620_o;
  /* helpers.vhdl:266:24  */
  assign n18622_o = n18617_o | n18621_o;
  /* helpers.vhdl:266:29  */
  assign n18623_o = n18565_o[19];
  /* helpers.vhdl:266:55  */
  assign n18624_o = n18565_o[18];
  /* helpers.vhdl:266:50  */
  assign n18625_o = ~n18624_o;
  /* helpers.vhdl:266:46  */
  assign n18626_o = n18623_o & n18625_o;
  /* helpers.vhdl:266:24  */
  assign n18627_o = n18622_o | n18626_o;
  /* helpers.vhdl:266:29  */
  assign n18628_o = n18565_o[21];
  /* helpers.vhdl:266:55  */
  assign n18629_o = n18565_o[20];
  /* helpers.vhdl:266:50  */
  assign n18630_o = ~n18629_o;
  /* helpers.vhdl:266:46  */
  assign n18631_o = n18628_o & n18630_o;
  /* helpers.vhdl:266:24  */
  assign n18632_o = n18627_o | n18631_o;
  /* helpers.vhdl:266:29  */
  assign n18633_o = n18565_o[23];
  /* helpers.vhdl:266:55  */
  assign n18634_o = n18565_o[22];
  /* helpers.vhdl:266:50  */
  assign n18635_o = ~n18634_o;
  /* helpers.vhdl:266:46  */
  assign n18636_o = n18633_o & n18635_o;
  /* helpers.vhdl:266:24  */
  assign n18637_o = n18632_o | n18636_o;
  /* helpers.vhdl:266:29  */
  assign n18638_o = n18565_o[25];
  /* helpers.vhdl:266:55  */
  assign n18639_o = n18565_o[24];
  /* helpers.vhdl:266:50  */
  assign n18640_o = ~n18639_o;
  /* helpers.vhdl:266:46  */
  assign n18641_o = n18638_o & n18640_o;
  /* helpers.vhdl:266:24  */
  assign n18642_o = n18637_o | n18641_o;
  /* helpers.vhdl:266:29  */
  assign n18643_o = n18565_o[27];
  /* helpers.vhdl:266:55  */
  assign n18644_o = n18565_o[26];
  /* helpers.vhdl:266:50  */
  assign n18645_o = ~n18644_o;
  /* helpers.vhdl:266:46  */
  assign n18646_o = n18643_o & n18645_o;
  /* helpers.vhdl:266:24  */
  assign n18647_o = n18642_o | n18646_o;
  /* helpers.vhdl:266:29  */
  assign n18648_o = n18565_o[29];
  /* helpers.vhdl:266:55  */
  assign n18649_o = n18565_o[28];
  /* helpers.vhdl:266:50  */
  assign n18650_o = ~n18649_o;
  /* helpers.vhdl:266:46  */
  assign n18651_o = n18648_o & n18650_o;
  /* helpers.vhdl:266:24  */
  assign n18652_o = n18647_o | n18651_o;
  /* helpers.vhdl:266:29  */
  assign n18653_o = n18565_o[31];
  /* helpers.vhdl:266:55  */
  assign n18654_o = n18565_o[30];
  /* helpers.vhdl:266:50  */
  assign n18655_o = ~n18654_o;
  /* helpers.vhdl:266:46  */
  assign n18656_o = n18653_o & n18655_o;
  /* helpers.vhdl:266:24  */
  assign n18657_o = n18652_o | n18656_o;
  /* helpers.vhdl:266:29  */
  assign n18658_o = n18565_o[33];
  /* helpers.vhdl:266:55  */
  assign n18659_o = n18565_o[32];
  /* helpers.vhdl:266:50  */
  assign n18660_o = ~n18659_o;
  /* helpers.vhdl:266:46  */
  assign n18661_o = n18658_o & n18660_o;
  /* helpers.vhdl:266:24  */
  assign n18662_o = n18657_o | n18661_o;
  /* helpers.vhdl:266:29  */
  assign n18663_o = n18565_o[35];
  /* helpers.vhdl:266:55  */
  assign n18664_o = n18565_o[34];
  /* helpers.vhdl:266:50  */
  assign n18665_o = ~n18664_o;
  /* helpers.vhdl:266:46  */
  assign n18666_o = n18663_o & n18665_o;
  /* helpers.vhdl:266:24  */
  assign n18667_o = n18662_o | n18666_o;
  /* helpers.vhdl:266:29  */
  assign n18668_o = n18565_o[37];
  /* helpers.vhdl:266:55  */
  assign n18669_o = n18565_o[36];
  /* helpers.vhdl:266:50  */
  assign n18670_o = ~n18669_o;
  /* helpers.vhdl:266:46  */
  assign n18671_o = n18668_o & n18670_o;
  /* helpers.vhdl:266:24  */
  assign n18672_o = n18667_o | n18671_o;
  /* helpers.vhdl:266:29  */
  assign n18673_o = n18565_o[39];
  /* helpers.vhdl:266:55  */
  assign n18674_o = n18565_o[38];
  /* helpers.vhdl:266:50  */
  assign n18675_o = ~n18674_o;
  /* helpers.vhdl:266:46  */
  assign n18676_o = n18673_o & n18675_o;
  /* helpers.vhdl:266:24  */
  assign n18677_o = n18672_o | n18676_o;
  /* helpers.vhdl:266:29  */
  assign n18678_o = n18565_o[41];
  /* helpers.vhdl:266:55  */
  assign n18679_o = n18565_o[40];
  /* helpers.vhdl:266:50  */
  assign n18680_o = ~n18679_o;
  /* helpers.vhdl:266:46  */
  assign n18681_o = n18678_o & n18680_o;
  /* helpers.vhdl:266:24  */
  assign n18682_o = n18677_o | n18681_o;
  /* helpers.vhdl:266:29  */
  assign n18683_o = n18565_o[43];
  /* helpers.vhdl:266:55  */
  assign n18684_o = n18565_o[42];
  /* helpers.vhdl:266:50  */
  assign n18685_o = ~n18684_o;
  /* helpers.vhdl:266:46  */
  assign n18686_o = n18683_o & n18685_o;
  /* helpers.vhdl:266:24  */
  assign n18687_o = n18682_o | n18686_o;
  /* helpers.vhdl:266:29  */
  assign n18688_o = n18565_o[45];
  /* helpers.vhdl:266:55  */
  assign n18689_o = n18565_o[44];
  /* helpers.vhdl:266:50  */
  assign n18690_o = ~n18689_o;
  /* helpers.vhdl:266:46  */
  assign n18691_o = n18688_o & n18690_o;
  /* helpers.vhdl:266:24  */
  assign n18692_o = n18687_o | n18691_o;
  /* helpers.vhdl:266:29  */
  assign n18693_o = n18565_o[47];
  /* helpers.vhdl:266:55  */
  assign n18694_o = n18565_o[46];
  /* helpers.vhdl:266:50  */
  assign n18695_o = ~n18694_o;
  /* helpers.vhdl:266:46  */
  assign n18696_o = n18693_o & n18695_o;
  /* helpers.vhdl:266:24  */
  assign n18697_o = n18692_o | n18696_o;
  /* helpers.vhdl:266:29  */
  assign n18698_o = n18565_o[49];
  /* helpers.vhdl:266:55  */
  assign n18699_o = n18565_o[48];
  /* helpers.vhdl:266:50  */
  assign n18700_o = ~n18699_o;
  /* helpers.vhdl:266:46  */
  assign n18701_o = n18698_o & n18700_o;
  /* helpers.vhdl:266:24  */
  assign n18702_o = n18697_o | n18701_o;
  /* helpers.vhdl:266:29  */
  assign n18703_o = n18565_o[51];
  /* helpers.vhdl:266:55  */
  assign n18704_o = n18565_o[50];
  /* helpers.vhdl:266:50  */
  assign n18705_o = ~n18704_o;
  /* helpers.vhdl:266:46  */
  assign n18706_o = n18703_o & n18705_o;
  /* helpers.vhdl:266:24  */
  assign n18707_o = n18702_o | n18706_o;
  /* helpers.vhdl:266:29  */
  assign n18708_o = n18565_o[53];
  /* helpers.vhdl:266:55  */
  assign n18709_o = n18565_o[52];
  /* helpers.vhdl:266:50  */
  assign n18710_o = ~n18709_o;
  /* helpers.vhdl:266:46  */
  assign n18711_o = n18708_o & n18710_o;
  /* helpers.vhdl:266:24  */
  assign n18712_o = n18707_o | n18711_o;
  /* helpers.vhdl:266:29  */
  assign n18713_o = n18565_o[55];
  /* helpers.vhdl:266:55  */
  assign n18714_o = n18565_o[54];
  /* helpers.vhdl:266:50  */
  assign n18715_o = ~n18714_o;
  /* helpers.vhdl:266:46  */
  assign n18716_o = n18713_o & n18715_o;
  /* helpers.vhdl:266:24  */
  assign n18717_o = n18712_o | n18716_o;
  /* helpers.vhdl:266:29  */
  assign n18718_o = n18565_o[57];
  /* helpers.vhdl:266:55  */
  assign n18719_o = n18565_o[56];
  /* helpers.vhdl:266:50  */
  assign n18720_o = ~n18719_o;
  /* helpers.vhdl:266:46  */
  assign n18721_o = n18718_o & n18720_o;
  /* helpers.vhdl:266:24  */
  assign n18722_o = n18717_o | n18721_o;
  /* helpers.vhdl:266:29  */
  assign n18723_o = n18565_o[59];
  /* helpers.vhdl:266:55  */
  assign n18724_o = n18565_o[58];
  /* helpers.vhdl:266:50  */
  assign n18725_o = ~n18724_o;
  /* helpers.vhdl:266:46  */
  assign n18726_o = n18723_o & n18725_o;
  /* helpers.vhdl:266:24  */
  assign n18727_o = n18722_o | n18726_o;
  /* helpers.vhdl:266:29  */
  assign n18728_o = n18565_o[61];
  /* helpers.vhdl:266:55  */
  assign n18729_o = n18565_o[60];
  /* helpers.vhdl:266:50  */
  assign n18730_o = ~n18729_o;
  /* helpers.vhdl:266:46  */
  assign n18731_o = n18728_o & n18730_o;
  /* helpers.vhdl:266:24  */
  assign n18732_o = n18727_o | n18731_o;
  /* helpers.vhdl:266:29  */
  assign n18733_o = n18565_o[63];
  /* helpers.vhdl:266:55  */
  assign n18734_o = n18565_o[62];
  /* helpers.vhdl:266:50  */
  assign n18735_o = ~n18734_o;
  /* helpers.vhdl:266:46  */
  assign n18736_o = n18733_o & n18735_o;
  /* helpers.vhdl:266:24  */
  assign n18737_o = n18732_o | n18736_o;
  /* helpers.vhdl:266:29  */
  assign n18740_o = n18565_o[3];
  /* helpers.vhdl:266:55  */
  assign n18741_o = n18565_o[1];
  /* helpers.vhdl:266:50  */
  assign n18742_o = ~n18741_o;
  /* helpers.vhdl:266:46  */
  assign n18743_o = n18740_o & n18742_o;
  /* helpers.vhdl:266:24  */
  assign n18745_o = 1'b0 | n18743_o;
  /* helpers.vhdl:266:29  */
  assign n18747_o = n18565_o[7];
  /* helpers.vhdl:266:55  */
  assign n18748_o = n18565_o[5];
  /* helpers.vhdl:266:50  */
  assign n18749_o = ~n18748_o;
  /* helpers.vhdl:266:46  */
  assign n18750_o = n18747_o & n18749_o;
  /* helpers.vhdl:266:24  */
  assign n18751_o = n18745_o | n18750_o;
  /* helpers.vhdl:266:29  */
  assign n18752_o = n18565_o[11];
  /* helpers.vhdl:266:55  */
  assign n18753_o = n18565_o[9];
  /* helpers.vhdl:266:50  */
  assign n18754_o = ~n18753_o;
  /* helpers.vhdl:266:46  */
  assign n18755_o = n18752_o & n18754_o;
  /* helpers.vhdl:266:24  */
  assign n18756_o = n18751_o | n18755_o;
  /* helpers.vhdl:266:29  */
  assign n18757_o = n18565_o[15];
  /* helpers.vhdl:266:55  */
  assign n18758_o = n18565_o[13];
  /* helpers.vhdl:266:50  */
  assign n18759_o = ~n18758_o;
  /* helpers.vhdl:266:46  */
  assign n18760_o = n18757_o & n18759_o;
  /* helpers.vhdl:266:24  */
  assign n18761_o = n18756_o | n18760_o;
  /* helpers.vhdl:266:29  */
  assign n18762_o = n18565_o[19];
  /* helpers.vhdl:266:55  */
  assign n18763_o = n18565_o[17];
  /* helpers.vhdl:266:50  */
  assign n18764_o = ~n18763_o;
  /* helpers.vhdl:266:46  */
  assign n18765_o = n18762_o & n18764_o;
  /* helpers.vhdl:266:24  */
  assign n18766_o = n18761_o | n18765_o;
  /* helpers.vhdl:266:29  */
  assign n18767_o = n18565_o[23];
  /* helpers.vhdl:266:55  */
  assign n18768_o = n18565_o[21];
  /* helpers.vhdl:266:50  */
  assign n18769_o = ~n18768_o;
  /* helpers.vhdl:266:46  */
  assign n18770_o = n18767_o & n18769_o;
  /* helpers.vhdl:266:24  */
  assign n18771_o = n18766_o | n18770_o;
  /* helpers.vhdl:266:29  */
  assign n18772_o = n18565_o[27];
  /* helpers.vhdl:266:55  */
  assign n18773_o = n18565_o[25];
  /* helpers.vhdl:266:50  */
  assign n18774_o = ~n18773_o;
  /* helpers.vhdl:266:46  */
  assign n18775_o = n18772_o & n18774_o;
  /* helpers.vhdl:266:24  */
  assign n18776_o = n18771_o | n18775_o;
  /* helpers.vhdl:266:29  */
  assign n18777_o = n18565_o[31];
  /* helpers.vhdl:266:55  */
  assign n18778_o = n18565_o[29];
  /* helpers.vhdl:266:50  */
  assign n18779_o = ~n18778_o;
  /* helpers.vhdl:266:46  */
  assign n18780_o = n18777_o & n18779_o;
  /* helpers.vhdl:266:24  */
  assign n18781_o = n18776_o | n18780_o;
  /* helpers.vhdl:266:29  */
  assign n18782_o = n18565_o[35];
  /* helpers.vhdl:266:55  */
  assign n18783_o = n18565_o[33];
  /* helpers.vhdl:266:50  */
  assign n18784_o = ~n18783_o;
  /* helpers.vhdl:266:46  */
  assign n18785_o = n18782_o & n18784_o;
  /* helpers.vhdl:266:24  */
  assign n18786_o = n18781_o | n18785_o;
  /* helpers.vhdl:266:29  */
  assign n18787_o = n18565_o[39];
  /* helpers.vhdl:266:55  */
  assign n18788_o = n18565_o[37];
  /* helpers.vhdl:266:50  */
  assign n18789_o = ~n18788_o;
  /* helpers.vhdl:266:46  */
  assign n18790_o = n18787_o & n18789_o;
  /* helpers.vhdl:266:24  */
  assign n18791_o = n18786_o | n18790_o;
  /* helpers.vhdl:266:29  */
  assign n18792_o = n18565_o[43];
  /* helpers.vhdl:266:55  */
  assign n18793_o = n18565_o[41];
  /* helpers.vhdl:266:50  */
  assign n18794_o = ~n18793_o;
  /* helpers.vhdl:266:46  */
  assign n18795_o = n18792_o & n18794_o;
  /* helpers.vhdl:266:24  */
  assign n18796_o = n18791_o | n18795_o;
  /* helpers.vhdl:266:29  */
  assign n18797_o = n18565_o[47];
  /* helpers.vhdl:266:55  */
  assign n18798_o = n18565_o[45];
  /* helpers.vhdl:266:50  */
  assign n18799_o = ~n18798_o;
  /* helpers.vhdl:266:46  */
  assign n18800_o = n18797_o & n18799_o;
  /* helpers.vhdl:266:24  */
  assign n18801_o = n18796_o | n18800_o;
  /* helpers.vhdl:266:29  */
  assign n18802_o = n18565_o[51];
  /* helpers.vhdl:266:55  */
  assign n18803_o = n18565_o[49];
  /* helpers.vhdl:266:50  */
  assign n18804_o = ~n18803_o;
  /* helpers.vhdl:266:46  */
  assign n18805_o = n18802_o & n18804_o;
  /* helpers.vhdl:266:24  */
  assign n18806_o = n18801_o | n18805_o;
  /* helpers.vhdl:266:29  */
  assign n18807_o = n18565_o[55];
  /* helpers.vhdl:266:55  */
  assign n18808_o = n18565_o[53];
  /* helpers.vhdl:266:50  */
  assign n18809_o = ~n18808_o;
  /* helpers.vhdl:266:46  */
  assign n18810_o = n18807_o & n18809_o;
  /* helpers.vhdl:266:24  */
  assign n18811_o = n18806_o | n18810_o;
  /* helpers.vhdl:266:29  */
  assign n18812_o = n18565_o[59];
  /* helpers.vhdl:266:55  */
  assign n18813_o = n18565_o[57];
  /* helpers.vhdl:266:50  */
  assign n18814_o = ~n18813_o;
  /* helpers.vhdl:266:46  */
  assign n18815_o = n18812_o & n18814_o;
  /* helpers.vhdl:266:24  */
  assign n18816_o = n18811_o | n18815_o;
  /* helpers.vhdl:266:29  */
  assign n18817_o = n18565_o[63];
  /* helpers.vhdl:266:55  */
  assign n18818_o = n18565_o[61];
  /* helpers.vhdl:266:50  */
  assign n18819_o = ~n18818_o;
  /* helpers.vhdl:266:46  */
  assign n18820_o = n18817_o & n18819_o;
  /* helpers.vhdl:266:24  */
  assign n18821_o = n18816_o | n18820_o;
  /* helpers.vhdl:266:29  */
  assign n18823_o = n18565_o[7];
  /* helpers.vhdl:266:55  */
  assign n18824_o = n18565_o[3];
  /* helpers.vhdl:266:50  */
  assign n18825_o = ~n18824_o;
  /* helpers.vhdl:266:46  */
  assign n18826_o = n18823_o & n18825_o;
  /* helpers.vhdl:266:24  */
  assign n18828_o = 1'b0 | n18826_o;
  /* helpers.vhdl:266:29  */
  assign n18830_o = n18565_o[15];
  /* helpers.vhdl:266:55  */
  assign n18831_o = n18565_o[11];
  /* helpers.vhdl:266:50  */
  assign n18832_o = ~n18831_o;
  /* helpers.vhdl:266:46  */
  assign n18833_o = n18830_o & n18832_o;
  /* helpers.vhdl:266:24  */
  assign n18834_o = n18828_o | n18833_o;
  /* helpers.vhdl:266:29  */
  assign n18835_o = n18565_o[23];
  /* helpers.vhdl:266:55  */
  assign n18836_o = n18565_o[19];
  /* helpers.vhdl:266:50  */
  assign n18837_o = ~n18836_o;
  /* helpers.vhdl:266:46  */
  assign n18838_o = n18835_o & n18837_o;
  /* helpers.vhdl:266:24  */
  assign n18839_o = n18834_o | n18838_o;
  /* helpers.vhdl:266:29  */
  assign n18840_o = n18565_o[31];
  /* helpers.vhdl:266:55  */
  assign n18841_o = n18565_o[27];
  /* helpers.vhdl:266:50  */
  assign n18842_o = ~n18841_o;
  /* helpers.vhdl:266:46  */
  assign n18843_o = n18840_o & n18842_o;
  /* helpers.vhdl:266:24  */
  assign n18844_o = n18839_o | n18843_o;
  /* helpers.vhdl:266:29  */
  assign n18845_o = n18565_o[39];
  /* helpers.vhdl:266:55  */
  assign n18846_o = n18565_o[35];
  /* helpers.vhdl:266:50  */
  assign n18847_o = ~n18846_o;
  /* helpers.vhdl:266:46  */
  assign n18848_o = n18845_o & n18847_o;
  /* helpers.vhdl:266:24  */
  assign n18849_o = n18844_o | n18848_o;
  /* helpers.vhdl:266:29  */
  assign n18850_o = n18565_o[47];
  /* helpers.vhdl:266:55  */
  assign n18851_o = n18565_o[43];
  /* helpers.vhdl:266:50  */
  assign n18852_o = ~n18851_o;
  /* helpers.vhdl:266:46  */
  assign n18853_o = n18850_o & n18852_o;
  /* helpers.vhdl:266:24  */
  assign n18854_o = n18849_o | n18853_o;
  /* helpers.vhdl:266:29  */
  assign n18855_o = n18565_o[55];
  /* helpers.vhdl:266:55  */
  assign n18856_o = n18565_o[51];
  /* helpers.vhdl:266:50  */
  assign n18857_o = ~n18856_o;
  /* helpers.vhdl:266:46  */
  assign n18858_o = n18855_o & n18857_o;
  /* helpers.vhdl:266:24  */
  assign n18859_o = n18854_o | n18858_o;
  /* helpers.vhdl:266:29  */
  assign n18860_o = n18565_o[63];
  /* helpers.vhdl:266:55  */
  assign n18861_o = n18565_o[59];
  /* helpers.vhdl:266:50  */
  assign n18862_o = ~n18861_o;
  /* helpers.vhdl:266:46  */
  assign n18863_o = n18860_o & n18862_o;
  /* helpers.vhdl:266:24  */
  assign n18864_o = n18859_o | n18863_o;
  /* helpers.vhdl:266:29  */
  assign n18866_o = n18565_o[15];
  /* helpers.vhdl:266:55  */
  assign n18867_o = n18565_o[7];
  /* helpers.vhdl:266:50  */
  assign n18868_o = ~n18867_o;
  /* helpers.vhdl:266:46  */
  assign n18869_o = n18866_o & n18868_o;
  /* helpers.vhdl:266:24  */
  assign n18871_o = 1'b0 | n18869_o;
  /* helpers.vhdl:266:29  */
  assign n18873_o = n18565_o[31];
  /* helpers.vhdl:266:55  */
  assign n18874_o = n18565_o[23];
  /* helpers.vhdl:266:50  */
  assign n18875_o = ~n18874_o;
  /* helpers.vhdl:266:46  */
  assign n18876_o = n18873_o & n18875_o;
  /* helpers.vhdl:266:24  */
  assign n18877_o = n18871_o | n18876_o;
  /* helpers.vhdl:266:29  */
  assign n18878_o = n18565_o[47];
  /* helpers.vhdl:266:55  */
  assign n18879_o = n18565_o[39];
  /* helpers.vhdl:266:50  */
  assign n18880_o = ~n18879_o;
  /* helpers.vhdl:266:46  */
  assign n18881_o = n18878_o & n18880_o;
  /* helpers.vhdl:266:24  */
  assign n18882_o = n18877_o | n18881_o;
  /* helpers.vhdl:266:29  */
  assign n18883_o = n18565_o[63];
  /* helpers.vhdl:266:55  */
  assign n18884_o = n18565_o[55];
  /* helpers.vhdl:266:50  */
  assign n18885_o = ~n18884_o;
  /* helpers.vhdl:266:46  */
  assign n18886_o = n18883_o & n18885_o;
  /* helpers.vhdl:266:24  */
  assign n18887_o = n18882_o | n18886_o;
  /* helpers.vhdl:266:29  */
  assign n18889_o = n18565_o[31];
  /* helpers.vhdl:266:55  */
  assign n18890_o = n18565_o[15];
  /* helpers.vhdl:266:50  */
  assign n18891_o = ~n18890_o;
  /* helpers.vhdl:266:46  */
  assign n18892_o = n18889_o & n18891_o;
  /* helpers.vhdl:266:24  */
  assign n18894_o = 1'b0 | n18892_o;
  /* helpers.vhdl:266:29  */
  assign n18896_o = n18565_o[63];
  /* helpers.vhdl:266:55  */
  assign n18897_o = n18565_o[47];
  /* helpers.vhdl:266:50  */
  assign n18898_o = ~n18897_o;
  /* helpers.vhdl:266:46  */
  assign n18899_o = n18896_o & n18898_o;
  /* helpers.vhdl:266:24  */
  assign n18900_o = n18894_o | n18899_o;
  /* helpers.vhdl:266:29  */
  assign n18902_o = n18565_o[63];
  /* helpers.vhdl:266:55  */
  assign n18903_o = n18565_o[31];
  /* helpers.vhdl:266:50  */
  assign n18904_o = ~n18903_o;
  /* helpers.vhdl:266:46  */
  assign n18905_o = n18902_o & n18904_o;
  /* helpers.vhdl:266:24  */
  assign n18907_o = 1'b0 | n18905_o;
  assign n18909_o = {n18907_o, n18900_o, n18887_o, n18864_o, n18821_o, n18737_o};
  /* helpers.vhdl:244:36  */
  assign n18920_o = n18563_o[1];
  /* helpers.vhdl:244:32  */
  assign n18921_o = |(n18920_o);
  /* helpers.vhdl:244:28  */
  assign n18923_o = 1'b0 | n18921_o;
  /* helpers.vhdl:244:36  */
  assign n18925_o = n18563_o[3];
  /* helpers.vhdl:244:32  */
  assign n18926_o = |(n18925_o);
  /* helpers.vhdl:244:28  */
  assign n18927_o = n18923_o | n18926_o;
  /* helpers.vhdl:244:36  */
  assign n18928_o = n18563_o[5];
  /* helpers.vhdl:244:32  */
  assign n18929_o = |(n18928_o);
  /* helpers.vhdl:244:28  */
  assign n18930_o = n18927_o | n18929_o;
  /* helpers.vhdl:244:36  */
  assign n18931_o = n18563_o[7];
  /* helpers.vhdl:244:32  */
  assign n18932_o = |(n18931_o);
  /* helpers.vhdl:244:28  */
  assign n18933_o = n18930_o | n18932_o;
  /* helpers.vhdl:244:36  */
  assign n18934_o = n18563_o[9];
  /* helpers.vhdl:244:32  */
  assign n18935_o = |(n18934_o);
  /* helpers.vhdl:244:28  */
  assign n18936_o = n18933_o | n18935_o;
  /* helpers.vhdl:244:36  */
  assign n18937_o = n18563_o[11];
  /* helpers.vhdl:244:32  */
  assign n18938_o = |(n18937_o);
  /* helpers.vhdl:244:28  */
  assign n18939_o = n18936_o | n18938_o;
  /* helpers.vhdl:244:36  */
  assign n18940_o = n18563_o[13];
  /* helpers.vhdl:244:32  */
  assign n18941_o = |(n18940_o);
  /* helpers.vhdl:244:28  */
  assign n18942_o = n18939_o | n18941_o;
  /* helpers.vhdl:244:36  */
  assign n18943_o = n18563_o[15];
  /* helpers.vhdl:244:32  */
  assign n18944_o = |(n18943_o);
  /* helpers.vhdl:244:28  */
  assign n18945_o = n18942_o | n18944_o;
  /* helpers.vhdl:244:36  */
  assign n18946_o = n18563_o[17];
  /* helpers.vhdl:244:32  */
  assign n18947_o = |(n18946_o);
  /* helpers.vhdl:244:28  */
  assign n18948_o = n18945_o | n18947_o;
  /* helpers.vhdl:244:36  */
  assign n18949_o = n18563_o[19];
  /* helpers.vhdl:244:32  */
  assign n18950_o = |(n18949_o);
  /* helpers.vhdl:244:28  */
  assign n18951_o = n18948_o | n18950_o;
  /* helpers.vhdl:244:36  */
  assign n18952_o = n18563_o[21];
  /* helpers.vhdl:244:32  */
  assign n18953_o = |(n18952_o);
  /* helpers.vhdl:244:28  */
  assign n18954_o = n18951_o | n18953_o;
  /* helpers.vhdl:244:36  */
  assign n18955_o = n18563_o[23];
  /* helpers.vhdl:244:32  */
  assign n18956_o = |(n18955_o);
  /* helpers.vhdl:244:28  */
  assign n18957_o = n18954_o | n18956_o;
  /* helpers.vhdl:244:36  */
  assign n18958_o = n18563_o[25];
  /* helpers.vhdl:244:32  */
  assign n18959_o = |(n18958_o);
  /* helpers.vhdl:244:28  */
  assign n18960_o = n18957_o | n18959_o;
  /* helpers.vhdl:244:36  */
  assign n18961_o = n18563_o[27];
  /* helpers.vhdl:244:32  */
  assign n18962_o = |(n18961_o);
  /* helpers.vhdl:244:28  */
  assign n18963_o = n18960_o | n18962_o;
  /* helpers.vhdl:244:36  */
  assign n18964_o = n18563_o[29];
  /* helpers.vhdl:244:32  */
  assign n18965_o = |(n18964_o);
  /* helpers.vhdl:244:28  */
  assign n18966_o = n18963_o | n18965_o;
  /* helpers.vhdl:244:36  */
  assign n18967_o = n18563_o[31];
  /* helpers.vhdl:244:32  */
  assign n18968_o = |(n18967_o);
  /* helpers.vhdl:244:28  */
  assign n18969_o = n18966_o | n18968_o;
  /* helpers.vhdl:244:36  */
  assign n18970_o = n18563_o[33];
  /* helpers.vhdl:244:32  */
  assign n18971_o = |(n18970_o);
  /* helpers.vhdl:244:28  */
  assign n18972_o = n18969_o | n18971_o;
  /* helpers.vhdl:244:36  */
  assign n18973_o = n18563_o[35];
  /* helpers.vhdl:244:32  */
  assign n18974_o = |(n18973_o);
  /* helpers.vhdl:244:28  */
  assign n18975_o = n18972_o | n18974_o;
  /* helpers.vhdl:244:36  */
  assign n18976_o = n18563_o[37];
  /* helpers.vhdl:244:32  */
  assign n18977_o = |(n18976_o);
  /* helpers.vhdl:244:28  */
  assign n18978_o = n18975_o | n18977_o;
  /* helpers.vhdl:244:36  */
  assign n18979_o = n18563_o[39];
  /* helpers.vhdl:244:32  */
  assign n18980_o = |(n18979_o);
  /* helpers.vhdl:244:28  */
  assign n18981_o = n18978_o | n18980_o;
  /* helpers.vhdl:244:36  */
  assign n18982_o = n18563_o[41];
  /* helpers.vhdl:244:32  */
  assign n18983_o = |(n18982_o);
  /* helpers.vhdl:244:28  */
  assign n18984_o = n18981_o | n18983_o;
  /* helpers.vhdl:244:36  */
  assign n18985_o = n18563_o[43];
  /* helpers.vhdl:244:32  */
  assign n18986_o = |(n18985_o);
  /* helpers.vhdl:244:28  */
  assign n18987_o = n18984_o | n18986_o;
  /* helpers.vhdl:244:36  */
  assign n18988_o = n18563_o[45];
  /* helpers.vhdl:244:32  */
  assign n18989_o = |(n18988_o);
  /* helpers.vhdl:244:28  */
  assign n18990_o = n18987_o | n18989_o;
  /* helpers.vhdl:244:36  */
  assign n18991_o = n18563_o[47];
  /* helpers.vhdl:244:32  */
  assign n18992_o = |(n18991_o);
  /* helpers.vhdl:244:28  */
  assign n18993_o = n18990_o | n18992_o;
  /* helpers.vhdl:244:36  */
  assign n18994_o = n18563_o[49];
  /* helpers.vhdl:244:32  */
  assign n18995_o = |(n18994_o);
  /* helpers.vhdl:244:28  */
  assign n18996_o = n18993_o | n18995_o;
  /* helpers.vhdl:244:36  */
  assign n18997_o = n18563_o[51];
  /* helpers.vhdl:244:32  */
  assign n18998_o = |(n18997_o);
  /* helpers.vhdl:244:28  */
  assign n18999_o = n18996_o | n18998_o;
  /* helpers.vhdl:244:36  */
  assign n19000_o = n18563_o[53];
  /* helpers.vhdl:244:32  */
  assign n19001_o = |(n19000_o);
  /* helpers.vhdl:244:28  */
  assign n19002_o = n18999_o | n19001_o;
  /* helpers.vhdl:244:36  */
  assign n19003_o = n18563_o[55];
  /* helpers.vhdl:244:32  */
  assign n19004_o = |(n19003_o);
  /* helpers.vhdl:244:28  */
  assign n19005_o = n19002_o | n19004_o;
  /* helpers.vhdl:244:36  */
  assign n19006_o = n18563_o[57];
  /* helpers.vhdl:244:32  */
  assign n19007_o = |(n19006_o);
  /* helpers.vhdl:244:28  */
  assign n19008_o = n19005_o | n19007_o;
  /* helpers.vhdl:244:36  */
  assign n19009_o = n18563_o[59];
  /* helpers.vhdl:244:32  */
  assign n19010_o = |(n19009_o);
  /* helpers.vhdl:244:28  */
  assign n19011_o = n19008_o | n19010_o;
  /* helpers.vhdl:244:36  */
  assign n19012_o = n18563_o[61];
  /* helpers.vhdl:244:32  */
  assign n19013_o = |(n19012_o);
  /* helpers.vhdl:244:28  */
  assign n19014_o = n19011_o | n19013_o;
  /* helpers.vhdl:244:36  */
  assign n19015_o = n18563_o[63];
  /* helpers.vhdl:244:32  */
  assign n19016_o = |(n19015_o);
  /* helpers.vhdl:244:28  */
  assign n19017_o = n19014_o | n19016_o;
  /* helpers.vhdl:244:36  */
  assign n19020_o = n18563_o[3:2];
  /* helpers.vhdl:244:32  */
  assign n19021_o = |(n19020_o);
  /* helpers.vhdl:244:28  */
  assign n19023_o = 1'b0 | n19021_o;
  /* helpers.vhdl:244:36  */
  assign n19025_o = n18563_o[7:6];
  /* helpers.vhdl:244:32  */
  assign n19026_o = |(n19025_o);
  /* helpers.vhdl:244:28  */
  assign n19027_o = n19023_o | n19026_o;
  /* helpers.vhdl:244:36  */
  assign n19028_o = n18563_o[11:10];
  /* helpers.vhdl:244:32  */
  assign n19029_o = |(n19028_o);
  /* helpers.vhdl:244:28  */
  assign n19030_o = n19027_o | n19029_o;
  /* helpers.vhdl:244:36  */
  assign n19031_o = n18563_o[15:14];
  /* helpers.vhdl:244:32  */
  assign n19032_o = |(n19031_o);
  /* helpers.vhdl:244:28  */
  assign n19033_o = n19030_o | n19032_o;
  /* helpers.vhdl:244:36  */
  assign n19034_o = n18563_o[19:18];
  /* helpers.vhdl:244:32  */
  assign n19035_o = |(n19034_o);
  /* helpers.vhdl:244:28  */
  assign n19036_o = n19033_o | n19035_o;
  /* helpers.vhdl:244:36  */
  assign n19037_o = n18563_o[23:22];
  /* helpers.vhdl:244:32  */
  assign n19038_o = |(n19037_o);
  /* helpers.vhdl:244:28  */
  assign n19039_o = n19036_o | n19038_o;
  /* helpers.vhdl:244:36  */
  assign n19040_o = n18563_o[27:26];
  /* helpers.vhdl:244:32  */
  assign n19041_o = |(n19040_o);
  /* helpers.vhdl:244:28  */
  assign n19042_o = n19039_o | n19041_o;
  /* helpers.vhdl:244:36  */
  assign n19043_o = n18563_o[31:30];
  /* helpers.vhdl:244:32  */
  assign n19044_o = |(n19043_o);
  /* helpers.vhdl:244:28  */
  assign n19045_o = n19042_o | n19044_o;
  /* helpers.vhdl:244:36  */
  assign n19046_o = n18563_o[35:34];
  /* helpers.vhdl:244:32  */
  assign n19047_o = |(n19046_o);
  /* helpers.vhdl:244:28  */
  assign n19048_o = n19045_o | n19047_o;
  /* helpers.vhdl:244:36  */
  assign n19049_o = n18563_o[39:38];
  /* helpers.vhdl:244:32  */
  assign n19050_o = |(n19049_o);
  /* helpers.vhdl:244:28  */
  assign n19051_o = n19048_o | n19050_o;
  /* helpers.vhdl:244:36  */
  assign n19052_o = n18563_o[43:42];
  /* helpers.vhdl:244:32  */
  assign n19053_o = |(n19052_o);
  /* helpers.vhdl:244:28  */
  assign n19054_o = n19051_o | n19053_o;
  /* helpers.vhdl:244:36  */
  assign n19055_o = n18563_o[47:46];
  /* helpers.vhdl:244:32  */
  assign n19056_o = |(n19055_o);
  /* helpers.vhdl:244:28  */
  assign n19057_o = n19054_o | n19056_o;
  /* helpers.vhdl:244:36  */
  assign n19058_o = n18563_o[51:50];
  /* helpers.vhdl:244:32  */
  assign n19059_o = |(n19058_o);
  /* helpers.vhdl:244:28  */
  assign n19060_o = n19057_o | n19059_o;
  /* helpers.vhdl:244:36  */
  assign n19061_o = n18563_o[55:54];
  /* helpers.vhdl:244:32  */
  assign n19062_o = |(n19061_o);
  /* helpers.vhdl:244:28  */
  assign n19063_o = n19060_o | n19062_o;
  /* helpers.vhdl:244:36  */
  assign n19064_o = n18563_o[59:58];
  /* helpers.vhdl:244:32  */
  assign n19065_o = |(n19064_o);
  /* helpers.vhdl:244:28  */
  assign n19066_o = n19063_o | n19065_o;
  /* helpers.vhdl:244:36  */
  assign n19067_o = n18563_o[63:62];
  /* helpers.vhdl:244:32  */
  assign n19068_o = |(n19067_o);
  /* helpers.vhdl:244:28  */
  assign n19069_o = n19066_o | n19068_o;
  /* helpers.vhdl:244:36  */
  assign n19071_o = n18563_o[7:4];
  /* helpers.vhdl:244:32  */
  assign n19072_o = |(n19071_o);
  /* helpers.vhdl:244:28  */
  assign n19074_o = 1'b0 | n19072_o;
  /* helpers.vhdl:244:36  */
  assign n19076_o = n18563_o[15:12];
  /* helpers.vhdl:244:32  */
  assign n19077_o = |(n19076_o);
  /* helpers.vhdl:244:28  */
  assign n19078_o = n19074_o | n19077_o;
  /* helpers.vhdl:244:36  */
  assign n19079_o = n18563_o[23:20];
  /* helpers.vhdl:244:32  */
  assign n19080_o = |(n19079_o);
  /* helpers.vhdl:244:28  */
  assign n19081_o = n19078_o | n19080_o;
  /* helpers.vhdl:244:36  */
  assign n19082_o = n18563_o[31:28];
  /* helpers.vhdl:244:32  */
  assign n19083_o = |(n19082_o);
  /* helpers.vhdl:244:28  */
  assign n19084_o = n19081_o | n19083_o;
  /* helpers.vhdl:244:36  */
  assign n19085_o = n18563_o[39:36];
  /* helpers.vhdl:244:32  */
  assign n19086_o = |(n19085_o);
  /* helpers.vhdl:244:28  */
  assign n19087_o = n19084_o | n19086_o;
  /* helpers.vhdl:244:36  */
  assign n19088_o = n18563_o[47:44];
  /* helpers.vhdl:244:32  */
  assign n19089_o = |(n19088_o);
  /* helpers.vhdl:244:28  */
  assign n19090_o = n19087_o | n19089_o;
  /* helpers.vhdl:244:36  */
  assign n19091_o = n18563_o[55:52];
  /* helpers.vhdl:244:32  */
  assign n19092_o = |(n19091_o);
  /* helpers.vhdl:244:28  */
  assign n19093_o = n19090_o | n19092_o;
  /* helpers.vhdl:244:36  */
  assign n19094_o = n18563_o[63:60];
  /* helpers.vhdl:244:32  */
  assign n19095_o = |(n19094_o);
  /* helpers.vhdl:244:28  */
  assign n19096_o = n19093_o | n19095_o;
  /* helpers.vhdl:244:36  */
  assign n19098_o = n18563_o[15:8];
  /* helpers.vhdl:244:32  */
  assign n19099_o = |(n19098_o);
  /* helpers.vhdl:244:28  */
  assign n19101_o = 1'b0 | n19099_o;
  /* helpers.vhdl:244:36  */
  assign n19103_o = n18563_o[31:24];
  /* helpers.vhdl:244:32  */
  assign n19104_o = |(n19103_o);
  /* helpers.vhdl:244:28  */
  assign n19105_o = n19101_o | n19104_o;
  /* helpers.vhdl:244:36  */
  assign n19106_o = n18563_o[47:40];
  /* helpers.vhdl:244:32  */
  assign n19107_o = |(n19106_o);
  /* helpers.vhdl:244:28  */
  assign n19108_o = n19105_o | n19107_o;
  /* helpers.vhdl:244:36  */
  assign n19109_o = n18563_o[63:56];
  /* helpers.vhdl:244:32  */
  assign n19110_o = |(n19109_o);
  /* helpers.vhdl:244:28  */
  assign n19111_o = n19108_o | n19110_o;
  /* helpers.vhdl:244:36  */
  assign n19113_o = n18563_o[31:16];
  /* helpers.vhdl:244:32  */
  assign n19114_o = |(n19113_o);
  /* helpers.vhdl:244:28  */
  assign n19116_o = 1'b0 | n19114_o;
  /* helpers.vhdl:244:36  */
  assign n19118_o = n18563_o[63:48];
  /* helpers.vhdl:244:32  */
  assign n19119_o = |(n19118_o);
  /* helpers.vhdl:244:28  */
  assign n19120_o = n19116_o | n19119_o;
  /* helpers.vhdl:244:36  */
  assign n19122_o = n18563_o[63:32];
  /* helpers.vhdl:244:32  */
  assign n19123_o = |(n19122_o);
  /* helpers.vhdl:244:28  */
  assign n19125_o = 1'b0 | n19123_o;
  assign n19127_o = {n19125_o, n19120_o, n19111_o, n19096_o, n19069_o, n19017_o};
  /* helpers.vhdl:287:19  */
  assign n19129_o = n18909_o[5:2];
  /* helpers.vhdl:287:38  */
  assign n19130_o = n19127_o[1:0];
  /* helpers.vhdl:287:32  */
  assign n19131_o = {n19129_o, n19130_o};
  assign n19134_o = n19131_o[0];
  /* fpu.vhdl:2522:13  */
  assign n19135_o = n17497_o ? 1'b1 : n19134_o;
  assign n19136_o = n19131_o[5:1];
  assign n19137_o = {n19136_o, n19135_o};
  /* fpu.vhdl:2526:42  */
  assign n19139_o = {1'b0, n19137_o};
  /* fpu.vhdl:2526:49  */
  assign n19141_o = n19139_o - 7'b0001001;
  /* fpu.vhdl:2526:24  */
  assign n19142_o = {{6{n19141_o[6]}}, n19141_o}; // sext
  /* fpu.vhdl:2520:9  */
  assign n19143_o = n17433_o ? n19142_o : n17174_o;
  /* fpu.vhdl:2529:14  */
  assign n19146_o = r[678];
  /* fpu.vhdl:2530:28  */
  assign n19147_o = r[462:399];
  /* fpu.vhdl:2532:36  */
  assign n19149_o = r[648];
  /* fpu.vhdl:2532:51  */
  assign n19150_o = r[650:649];
  /* fpu.vhdl:2532:67  */
  assign n19151_o = r[663:651];
  /* fpu.vhdl:2532:81  */
  assign n19152_o = r[462:399];
  /* fpu.vhdl:2533:36  */
  assign n19153_o = r[126];
  /* fpu.vhdl:2533:51  */
  assign n19154_o = r[697];
  /* fpu.vhdl:457:13  */
  assign n19163_o = n19150_o == 2'b00;
  /* fpu.vhdl:459:28  */
  assign n19164_o = n19152_o[54];
  /* fpu.vhdl:461:63  */
  assign n19165_o = n19151_o[10:0];  // trunc
  /* fpu.vhdl:461:79  */
  assign n19167_o = n19165_o + 11'b01111111111;
  assign n19168_o = n19160_o[62:52];
  /* fpu.vhdl:459:17  */
  assign n19169_o = n19164_o ? n19167_o : n19168_o;
  /* fpu.vhdl:463:49  */
  assign n19170_o = n19152_o[53:31];
  /* fpu.vhdl:464:32  */
  assign n19171_o = ~n19153_o;
  /* fpu.vhdl:465:52  */
  assign n19172_o = n19152_o[30:2];
  assign n19173_o = n19160_o[28:0];
  /* fpu.vhdl:464:17  */
  assign n19174_o = n19171_o ? n19172_o : n19173_o;
  /* fpu.vhdl:458:13  */
  assign n19176_o = n19150_o == 2'b01;
  /* fpu.vhdl:467:13  */
  assign n19179_o = n19150_o == 2'b10;
  /* fpu.vhdl:471:54  */
  assign n19181_o = n19152_o[53];
  /* fpu.vhdl:471:43  */
  assign n19182_o = n19154_o | n19181_o;
  /* fpu.vhdl:472:49  */
  assign n19183_o = n19152_o[52:31];
  /* fpu.vhdl:473:32  */
  assign n19184_o = ~n19153_o;
  /* fpu.vhdl:474:52  */
  assign n19185_o = n19152_o[30:2];
  assign n19186_o = n19160_o[28:0];
  /* fpu.vhdl:473:17  */
  assign n19187_o = n19184_o ? n19185_o : n19186_o;
  /* fpu.vhdl:469:13  */
  assign n19189_o = n19150_o == 2'b11;
  assign n19190_o = {n19189_o, n19179_o, n19176_o, n19163_o};
  assign n19191_o = n19160_o[28:0];
  /* fpu.vhdl:456:9  */
  always @*
    case (n19190_o)
      4'b1000: n19193_o = n19187_o;
      4'b0100: n19193_o = n19191_o;
      4'b0010: n19193_o = n19174_o;
      4'b0001: n19193_o = n19191_o;
      default: n19193_o = 29'bX;
    endcase
  assign n19194_o = n19170_o[21:0];
  assign n19195_o = n19160_o[50:29];
  /* fpu.vhdl:456:9  */
  always @*
    case (n19190_o)
      4'b1000: n19197_o = n19183_o;
      4'b0100: n19197_o = n19195_o;
      4'b0010: n19197_o = n19194_o;
      4'b0001: n19197_o = n19195_o;
      default: n19197_o = 22'bX;
    endcase
  assign n19198_o = n19170_o[22];
  assign n19199_o = n19160_o[51];
  /* fpu.vhdl:456:9  */
  always @*
    case (n19190_o)
      4'b1000: n19201_o = n19182_o;
      4'b0100: n19201_o = n19199_o;
      4'b0010: n19201_o = n19198_o;
      4'b0001: n19201_o = n19199_o;
      default: n19201_o = 1'bX;
    endcase
  assign n19202_o = n19160_o[62:52];
  /* fpu.vhdl:456:9  */
  always @*
    case (n19190_o)
      4'b1000: n19204_o = 11'b11111111111;
      4'b0100: n19204_o = 11'b11111111111;
      4'b0010: n19204_o = n19169_o;
      4'b0001: n19204_o = n19202_o;
      default: n19204_o = 11'bX;
    endcase
  assign n19208_o = {n19149_o, n19204_o, n19201_o, n19197_o, n19193_o};
  /* fpu.vhdl:2529:9  */
  assign n19209_o = n19146_o ? n19147_o : n19208_o;
  /* fpu.vhdl:2535:14  */
  assign n19210_o = r[696];
  /* fpu.vhdl:2536:64  */
  assign n19212_o = r[648];
  /* fpu.vhdl:2536:79  */
  assign n19213_o = r[650:649];
  /* fpu.vhdl:2537:65  */
  assign n19214_o = r[453];
  /* fpu.vhdl:2537:80  */
  assign n19215_o = r[699];
  /* fpu.vhdl:2537:74  */
  assign n19216_o = ~n19215_o;
  /* fpu.vhdl:2537:70  */
  assign n19217_o = n19214_o & n19216_o;
  /* fpu.vhdl:524:29  */
  assign n19223_o = {n19212_o, 4'b0010};
  /* fpu.vhdl:523:13  */
  assign n19225_o = n19213_o == 2'b00;
  /* fpu.vhdl:526:25  */
  assign n19226_o = ~n19217_o;
  /* fpu.vhdl:526:38  */
  assign n19227_o = {n19226_o, n19212_o};
  /* fpu.vhdl:526:48  */
  assign n19228_o = ~n19212_o;
  /* fpu.vhdl:526:45  */
  assign n19229_o = {n19227_o, n19228_o};
  /* fpu.vhdl:526:58  */
  assign n19231_o = {n19229_o, 2'b00};
  /* fpu.vhdl:525:13  */
  assign n19233_o = n19213_o == 2'b01;
  /* fpu.vhdl:528:28  */
  assign n19235_o = {1'b0, n19212_o};
  /* fpu.vhdl:528:38  */
  assign n19236_o = ~n19212_o;
  /* fpu.vhdl:528:35  */
  assign n19237_o = {n19235_o, n19236_o};
  /* fpu.vhdl:528:48  */
  assign n19239_o = {n19237_o, 2'b01};
  /* fpu.vhdl:527:13  */
  assign n19241_o = n19213_o == 2'b10;
  /* fpu.vhdl:529:13  */
  assign n19244_o = n19213_o == 2'b11;
  assign n19245_o = {n19244_o, n19241_o, n19233_o, n19225_o};
  /* fpu.vhdl:522:9  */
  always @*
    case (n19245_o)
      4'b1000: n19247_o = 5'b10001;
      4'b0100: n19247_o = n19239_o;
      4'b0010: n19247_o = n19231_o;
      4'b0001: n19247_o = n19223_o;
      default: n19247_o = 5'bX;
    endcase
  assign n19248_o = {n17056_o, n17050_o, n17042_o, n17034_o, n17026_o};
  /* fpu.vhdl:2535:9  */
  assign n19249_o = n19210_o ? n19247_o : n19248_o;
  assign n19250_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, n17538_o, n17204_o, n13473_o, n17202_o, n17196_o, n17190_o, n17184_o, n17178_o, n17537_o, n19143_o, n18406_o, n17519_o, n17644_o, n17651_o, n18373_o, result, n18400_o, n18403_o, n18389_o, n18395_o, n18378_o, n18384_o, n17154_o, n17148_o, n17142_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n19249_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n13556_o, n17542_o, 1'b0, n17541_o};
  /* fpu.vhdl:2540:42  */
  assign n19251_o = n19250_o[151:146];
  /* fpu.vhdl:2540:31  */
  assign n19252_o = |(n19251_o);
  assign n19253_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, n17538_o, n17204_o, n13473_o, n17202_o, n17196_o, n17190_o, n17184_o, n17178_o, n17537_o, n19143_o, n18406_o, n17519_o, n17644_o, n17651_o, n18373_o, result, n18400_o, n18403_o, n18389_o, n18395_o, n18378_o, n18384_o, n17154_o, n17148_o, n17142_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n19249_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n13556_o, n17542_o, 1'b0, n17541_o};
  /* fpu.vhdl:2541:42  */
  assign n19254_o = n19253_o[137:135];
  /* fpu.vhdl:2541:31  */
  assign n19255_o = |(n19254_o);
  /* fpu.vhdl:2540:77  */
  assign n19256_o = n19252_o | n19255_o;
  assign n19257_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, n17538_o, n17204_o, n13473_o, n17202_o, n17196_o, n17190_o, n17184_o, n17178_o, n17537_o, n19143_o, n18406_o, n17519_o, n17644_o, n17651_o, n18373_o, result, n18400_o, n18403_o, n18389_o, n18395_o, n18378_o, n18384_o, n17154_o, n17148_o, n19256_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n19249_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n13556_o, n17542_o, 1'b0, n17541_o};
  /* fpu.vhdl:2542:42  */
  assign n19258_o = n19257_o[156:152];
  assign n19259_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, n17538_o, n17204_o, n13473_o, n17202_o, n17196_o, n17190_o, n17184_o, n17178_o, n17537_o, n19143_o, n18406_o, n17519_o, n17644_o, n17651_o, n18373_o, result, n18400_o, n18403_o, n18389_o, n18395_o, n18378_o, n18384_o, n17154_o, n17148_o, n19256_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n19249_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n13556_o, n17542_o, 1'b0, n17541_o};
  /* fpu.vhdl:2543:42  */
  assign n19260_o = n19259_o[134:130];
  /* fpu.vhdl:2542:69  */
  assign n19261_o = n19258_o & n19260_o;
  /* fpu.vhdl:2542:31  */
  assign n19262_o = |(n19261_o);
  assign n19263_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, n17538_o, n17204_o, n13473_o, n17202_o, n17196_o, n17190_o, n17184_o, n17178_o, n17537_o, n19143_o, n18406_o, n17519_o, n17644_o, n17651_o, n18373_o, result, n18400_o, n18403_o, n18389_o, n18395_o, n18378_o, n18384_o, n17154_o, n19262_o, n19256_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n19249_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n13556_o, n17542_o, 1'b0, n17541_o};
  /* fpu.vhdl:2545:21  */
  assign n19264_o = n19263_o[156:152];
  /* fpu.vhdl:2545:58  */
  assign n19265_o = r[695:691];
  /* fpu.vhdl:2545:52  */
  assign n19266_o = ~n19265_o;
  /* fpu.vhdl:2545:48  */
  assign n19267_o = n19264_o & n19266_o;
  /* fpu.vhdl:2545:67  */
  assign n19269_o = n19267_o != 5'b00000;
  /* fpu.vhdl:2544:28  */
  assign n19270_o = n17546_o & n19269_o;
  /* fpu.vhdl:2544:9  */
  assign n19272_o = n19270_o ? 1'b1 : n17154_o;
  /* fpu.vhdl:2548:14  */
  assign n19273_o = r[124];
  assign n19274_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, n17538_o, n17204_o, n13473_o, n17202_o, n17196_o, n17190_o, n17184_o, n17178_o, n17537_o, n19143_o, n18406_o, n17519_o, n17644_o, n17651_o, n18373_o, result, n18400_o, n18403_o, n18389_o, n18395_o, n18378_o, n18384_o, n19272_o, n19262_o, n19256_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n19249_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n13556_o, n17542_o, 1'b0, n17541_o};
  /* fpu.vhdl:2549:35  */
  assign n19275_o = n19274_o[158:155];
  assign n19276_o = {n17202_o, n17196_o, n17190_o, n17184_o};
  /* fpu.vhdl:2548:9  */
  assign n19277_o = n19273_o ? n19275_o : n19276_o;
  assign n19278_o = r[9];
  assign n19284_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, n17538_o, n17204_o, n13473_o, n19277_o, n17178_o, n17537_o, n19143_o, n18406_o, n17519_o, n17644_o, n17651_o, n18373_o, result, n18400_o, n18403_o, n18389_o, n18395_o, n18378_o, n18384_o, n19272_o, n19262_o, n19256_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n19249_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n17393_o, n19278_o, n17542_o, 1'b0, n17541_o};
  /* fpu.vhdl:2560:28  */
  assign n19285_o = n19284_o[8];
  assign n19286_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, n17538_o, n17204_o, n13473_o, n19277_o, n17178_o, n17537_o, n19143_o, n18406_o, n17519_o, n17644_o, n17651_o, n18373_o, result, n18400_o, n18403_o, n18389_o, n18395_o, n18378_o, n18384_o, n19272_o, n19262_o, n19256_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n19249_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n17393_o, n19278_o, n17542_o, 1'b0, n17541_o};
  /* fpu.vhdl:2560:50  */
  assign n19287_o = n19286_o[157];
  /* fpu.vhdl:2560:39  */
  assign n19288_o = n19285_o & n19287_o;
  /* fpu.vhdl:2560:68  */
  assign n19289_o = r[123];
  /* fpu.vhdl:2560:62  */
  assign n19290_o = n19288_o & n19289_o;
  assign n19291_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, n17538_o, n17204_o, n13473_o, n19277_o, n17178_o, n17537_o, n19143_o, n18406_o, n17519_o, n17644_o, n17651_o, n18373_o, result, n18400_o, n18403_o, n18389_o, n18395_o, n18378_o, n18384_o, n19272_o, n19262_o, n19256_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n19249_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n17393_o, n19290_o, n17542_o, 1'b0, n17541_o};
  /* fpu.vhdl:2561:18  */
  assign n19292_o = n19291_o[6:0];
  /* fpu.vhdl:2561:24  */
  assign n19294_o = n19292_o != 7'b0000000;
  assign n19295_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, n17538_o, n17204_o, n13473_o, n19277_o, n17178_o, n17537_o, n19143_o, n18406_o, n17519_o, n17644_o, n17651_o, n18373_o, result, n18400_o, n18403_o, n18389_o, n18395_o, n18378_o, n18384_o, n19272_o, n19262_o, n19256_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n19249_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n17393_o, n19290_o, n17542_o, 1'b0, n17541_o};
  /* fpu.vhdl:2561:37  */
  assign n19296_o = n19295_o[9];
  /* fpu.vhdl:2561:32  */
  assign n19297_o = n19294_o | n19296_o;
  /* fpu.vhdl:2561:13  */
  assign n19299_o = n19297_o ? 1'b1 : 1'b0;
  assign n19300_o = {1'b1, 1'b0, 1'b0, 7'b0000000};
  assign n19301_o = n19300_o[6:0];
  /* fpu.vhdl:2553:9  */
  assign n19302_o = n17393_o ? n19301_o : n17541_o;
  assign n19303_o = n19300_o[7];
  /* fpu.vhdl:2553:9  */
  assign n19304_o = n17393_o ? n19303_o : n19299_o;
  assign n19305_o = n19300_o[8];
  /* fpu.vhdl:2553:9  */
  assign n19306_o = n17393_o ? n19305_o : n17542_o;
  assign n19307_o = n19300_o[9];
  /* fpu.vhdl:2553:9  */
  assign n19308_o = n17393_o ? n19307_o : n19290_o;
  /* fpu.vhdl:2553:9  */
  assign n19309_o = n17393_o ? 1'b0 : n17537_o;
  assign n19310_o = {n17280_o, n17278_o, n17525_o, n17272_o, n17269_o, n17266_o, n17263_o, n17261_o, n17259_o, n17255_o, n17251_o, n17245_o, n17239_o, n17234_o, n17340_o, n17229_o, n17224_o, n17219_o, n17214_o, n17209_o, n17538_o, n17204_o, n13473_o, n19277_o, n17178_o, n19309_o, n19143_o, n18406_o, n17519_o, n17644_o, n17651_o, n18373_o, result, n18400_o, n18403_o, n18389_o, n18395_o, n18378_o, n18384_o, n19272_o, n19262_o, n19256_o, n17136_o, n17130_o, n17509_o, n17118_o, n17112_o, n17106_o, n17100_o, n17093_o, n17086_o, n17080_o, n17074_o, n17065_o, n19249_o, n17018_o, n17012_o, n17006_o, n17000_o, n16994_o, n16987_o, n16980_o, n16973_o, n16966_o, n16959_o, n16953_o, n16946_o, n13467_o, n17393_o, n19308_o, n19306_o, n19304_o, n19302_o};
  /* fpu.vhdl:544:9  */
  always @(posedge clk)
    n19318_q <= n13017_o;
  assign n19320_o = {msel_inv, 1'b0, n17641_o, n17585_o, n17564_o, n16885_o};
  /* fpu.vhdl:564:9  */
  always @(posedge clk)
    n19321_q <= n13037_o;
  /* fpu.vhdl:564:9  */
  assign n19322_o = {n13043_o, n13042_o};
  assign n19323_o = {n13096_o, n13074_o, 12'b011100000000, n13071_o, n13056_o, n13055_o, fp_result, n13050_o, n13049_o, n13048_o, n13072_o, n13047_o};
  reg [17:0] n19324[1023:0] ; // memory
  initial begin
    n19324[1023] = 18'b111111110000000001;
    n19324[1022] = 18'b111111010000010001;
    n19324[1021] = 18'b111110110000110001;
    n19324[1020] = 18'b111110010001100000;
    n19324[1019] = 18'b111101110010011111;
    n19324[1018] = 18'b111101010011101100;
    n19324[1017] = 18'b111100110101001001;
    n19324[1016] = 18'b111100010110110101;
    n19324[1015] = 18'b111011111000101111;
    n19324[1014] = 18'b111011011010111000;
    n19324[1013] = 18'b111010111101001111;
    n19324[1012] = 18'b111010011111110100;
    n19324[1011] = 18'b111010000010100111;
    n19324[1010] = 18'b111001100101101000;
    n19324[1009] = 18'b111001001000110111;
    n19324[1008] = 18'b111000101100010100;
    n19324[1007] = 18'b111000001111111110;
    n19324[1006] = 18'b110111110011110101;
    n19324[1005] = 18'b110111010111111001;
    n19324[1004] = 18'b110110111100001010;
    n19324[1003] = 18'b110110100000101000;
    n19324[1002] = 18'b110110000101010011;
    n19324[1001] = 18'b110101101010001010;
    n19324[1000] = 18'b110101001111001110;
    n19324[999] = 18'b110100110100011110;
    n19324[998] = 18'b110100011001111010;
    n19324[997] = 18'b110011111111100011;
    n19324[996] = 18'b110011100101010111;
    n19324[995] = 18'b110011001011010111;
    n19324[994] = 18'b110010110001100010;
    n19324[993] = 18'b110010010111111001;
    n19324[992] = 18'b110001111110011100;
    n19324[991] = 18'b110001100101001010;
    n19324[990] = 18'b110001001100000011;
    n19324[989] = 18'b110000110011000111;
    n19324[988] = 18'b110000011010010110;
    n19324[987] = 18'b110000000001110000;
    n19324[986] = 18'b101111101001010100;
    n19324[985] = 18'b101111010001000011;
    n19324[984] = 18'b101110111000111101;
    n19324[983] = 18'b101110100001000001;
    n19324[982] = 18'b101110001001010000;
    n19324[981] = 18'b101101110001101000;
    n19324[980] = 18'b101101011010001011;
    n19324[979] = 18'b101101000010111000;
    n19324[978] = 18'b101100101011101110;
    n19324[977] = 18'b101100010100101110;
    n19324[976] = 18'b101011111101111001;
    n19324[975] = 18'b101011100111001100;
    n19324[974] = 18'b101011010000101001;
    n19324[973] = 18'b101010111010010000;
    n19324[972] = 18'b101010100100000000;
    n19324[971] = 18'b101010001101111001;
    n19324[970] = 18'b101001110111111011;
    n19324[969] = 18'b101001100010000111;
    n19324[968] = 18'b101001001100011011;
    n19324[967] = 18'b101000110110111000;
    n19324[966] = 18'b101000100001011110;
    n19324[965] = 18'b101000001100001101;
    n19324[964] = 18'b100111110111000100;
    n19324[963] = 18'b100111100010000100;
    n19324[962] = 18'b100111001101001101;
    n19324[961] = 18'b100110111000011101;
    n19324[960] = 18'b100110100011110110;
    n19324[959] = 18'b100110001111011000;
    n19324[958] = 18'b100101111011000001;
    n19324[957] = 18'b100101100110110011;
    n19324[956] = 18'b100101010010101100;
    n19324[955] = 18'b100100111110101101;
    n19324[954] = 18'b100100101010110111;
    n19324[953] = 18'b100100010111001000;
    n19324[952] = 18'b100100000011100001;
    n19324[951] = 18'b100011110000000001;
    n19324[950] = 18'b100011011100101001;
    n19324[949] = 18'b100011001001011001;
    n19324[948] = 18'b100010110110010000;
    n19324[947] = 18'b100010100011001110;
    n19324[946] = 18'b100010010000010011;
    n19324[945] = 18'b100001111101100000;
    n19324[944] = 18'b100001101010110100;
    n19324[943] = 18'b100001011000001111;
    n19324[942] = 18'b100001000101110010;
    n19324[941] = 18'b100000110011011011;
    n19324[940] = 18'b100000100001001011;
    n19324[939] = 18'b100000001111000010;
    n19324[938] = 18'b011111111101000000;
    n19324[937] = 18'b011111101011000100;
    n19324[936] = 18'b011111011001001111;
    n19324[935] = 18'b011111000111100001;
    n19324[934] = 18'b011110110101111001;
    n19324[933] = 18'b011110100100011000;
    n19324[932] = 18'b011110010010111110;
    n19324[931] = 18'b011110000001101001;
    n19324[930] = 18'b011101110000011011;
    n19324[929] = 18'b011101011111010100;
    n19324[928] = 18'b011101001110010010;
    n19324[927] = 18'b011100111101010111;
    n19324[926] = 18'b011100101100100010;
    n19324[925] = 18'b011100011011110011;
    n19324[924] = 18'b011100001011001010;
    n19324[923] = 18'b011011111010100111;
    n19324[922] = 18'b011011101010001010;
    n19324[921] = 18'b011011011001110010;
    n19324[920] = 18'b011011001001100001;
    n19324[919] = 18'b011010111001010101;
    n19324[918] = 18'b011010101001010000;
    n19324[917] = 18'b011010011001001111;
    n19324[916] = 18'b011010001001010101;
    n19324[915] = 18'b011001111001100000;
    n19324[914] = 18'b011001101001110000;
    n19324[913] = 18'b011001011010000110;
    n19324[912] = 18'b011001001010100010;
    n19324[911] = 18'b011000111011000011;
    n19324[910] = 18'b011000101011101001;
    n19324[909] = 18'b011000011100010101;
    n19324[908] = 18'b011000001101000101;
    n19324[907] = 18'b010111111101111100;
    n19324[906] = 18'b010111101110110111;
    n19324[905] = 18'b010111011111110111;
    n19324[904] = 18'b010111010000111101;
    n19324[903] = 18'b010111000010000111;
    n19324[902] = 18'b010110110011010111;
    n19324[901] = 18'b010110100100101100;
    n19324[900] = 18'b010110010110000101;
    n19324[899] = 18'b010110000111100100;
    n19324[898] = 18'b010101111001000111;
    n19324[897] = 18'b010101101010110000;
    n19324[896] = 18'b010101011100011101;
    n19324[895] = 18'b010101001110001110;
    n19324[894] = 18'b010101000000000101;
    n19324[893] = 18'b010100110010000000;
    n19324[892] = 18'b010100100100000000;
    n19324[891] = 18'b010100010110000100;
    n19324[890] = 18'b010100001000001101;
    n19324[889] = 18'b010011111010011011;
    n19324[888] = 18'b010011101100101101;
    n19324[887] = 18'b010011011111000011;
    n19324[886] = 18'b010011010001011110;
    n19324[885] = 18'b010011000011111110;
    n19324[884] = 18'b010010110110100010;
    n19324[883] = 18'b010010101001001010;
    n19324[882] = 18'b010010011011110110;
    n19324[881] = 18'b010010001110100111;
    n19324[880] = 18'b010010000001011100;
    n19324[879] = 18'b010001110100010101;
    n19324[878] = 18'b010001100111010010;
    n19324[877] = 18'b010001011010010100;
    n19324[876] = 18'b010001001101011001;
    n19324[875] = 18'b010001000000100011;
    n19324[874] = 18'b010000110011110001;
    n19324[873] = 18'b010000100111000010;
    n19324[872] = 18'b010000011010011000;
    n19324[871] = 18'b010000001101110010;
    n19324[870] = 18'b010000000001010000;
    n19324[869] = 18'b001111110100110001;
    n19324[868] = 18'b001111101000010111;
    n19324[867] = 18'b001111011100000000;
    n19324[866] = 18'b001111001111101101;
    n19324[865] = 18'b001111000011011110;
    n19324[864] = 18'b001110110111010011;
    n19324[863] = 18'b001110101011001011;
    n19324[862] = 18'b001110011111000111;
    n19324[861] = 18'b001110010011000111;
    n19324[860] = 18'b001110000111001010;
    n19324[859] = 18'b001101111011010010;
    n19324[858] = 18'b001101101111011100;
    n19324[857] = 18'b001101100011101011;
    n19324[856] = 18'b001101010111111100;
    n19324[855] = 18'b001101001100010010;
    n19324[854] = 18'b001101000000101011;
    n19324[853] = 18'b001100110101000111;
    n19324[852] = 18'b001100101001100111;
    n19324[851] = 18'b001100011110001010;
    n19324[850] = 18'b001100010010110001;
    n19324[849] = 18'b001100000111011011;
    n19324[848] = 18'b001011111100001001;
    n19324[847] = 18'b001011110000111010;
    n19324[846] = 18'b001011100101101110;
    n19324[845] = 18'b001011011010100101;
    n19324[844] = 18'b001011001111100000;
    n19324[843] = 18'b001011000100011110;
    n19324[842] = 18'b001010111001011111;
    n19324[841] = 18'b001010101110100011;
    n19324[840] = 18'b001010100011101011;
    n19324[839] = 18'b001010011000110110;
    n19324[838] = 18'b001010001110000011;
    n19324[837] = 18'b001010000011010100;
    n19324[836] = 18'b001001111000101000;
    n19324[835] = 18'b001001101110000000;
    n19324[834] = 18'b001001100011011010;
    n19324[833] = 18'b001001011000110111;
    n19324[832] = 18'b001001001110010111;
    n19324[831] = 18'b001001000011111011;
    n19324[830] = 18'b001000111001100001;
    n19324[829] = 18'b001000101111001010;
    n19324[828] = 18'b001000100100110110;
    n19324[827] = 18'b001000011010100101;
    n19324[826] = 18'b001000010000010111;
    n19324[825] = 18'b001000000110001100;
    n19324[824] = 18'b000111111100000100;
    n19324[823] = 18'b000111110001111110;
    n19324[822] = 18'b000111100111111100;
    n19324[821] = 18'b000111011101111100;
    n19324[820] = 18'b000111010011111111;
    n19324[819] = 18'b000111001010000100;
    n19324[818] = 18'b000111000000001101;
    n19324[817] = 18'b000110110110011000;
    n19324[816] = 18'b000110101100100110;
    n19324[815] = 18'b000110100010110110;
    n19324[814] = 18'b000110011001001010;
    n19324[813] = 18'b000110001111100000;
    n19324[812] = 18'b000110000101111000;
    n19324[811] = 18'b000101111100010011;
    n19324[810] = 18'b000101110010110001;
    n19324[809] = 18'b000101101001010010;
    n19324[808] = 18'b000101011111110101;
    n19324[807] = 18'b000101010110011010;
    n19324[806] = 18'b000101001101000010;
    n19324[805] = 18'b000101000011101101;
    n19324[804] = 18'b000100111010011010;
    n19324[803] = 18'b000100110001001010;
    n19324[802] = 18'b000100100111111100;
    n19324[801] = 18'b000100011110110000;
    n19324[800] = 18'b000100010101100111;
    n19324[799] = 18'b000100001100100001;
    n19324[798] = 18'b000100000011011101;
    n19324[797] = 18'b000011111010011011;
    n19324[796] = 18'b000011110001011100;
    n19324[795] = 18'b000011101000011111;
    n19324[794] = 18'b000011011111100100;
    n19324[793] = 18'b000011010110101100;
    n19324[792] = 18'b000011001101110110;
    n19324[791] = 18'b000011000101000010;
    n19324[790] = 18'b000010111100010001;
    n19324[789] = 18'b000010110011100010;
    n19324[788] = 18'b000010101010110101;
    n19324[787] = 18'b000010100010001011;
    n19324[786] = 18'b000010011001100011;
    n19324[785] = 18'b000010010000111101;
    n19324[784] = 18'b000010001000011001;
    n19324[783] = 18'b000001111111110111;
    n19324[782] = 18'b000001110111011000;
    n19324[781] = 18'b000001101110111011;
    n19324[780] = 18'b000001100110100000;
    n19324[779] = 18'b000001011110000111;
    n19324[778] = 18'b000001010101110000;
    n19324[777] = 18'b000001001101011011;
    n19324[776] = 18'b000001000101001001;
    n19324[775] = 18'b000000111100111001;
    n19324[774] = 18'b000000110100101010;
    n19324[773] = 18'b000000101100011110;
    n19324[772] = 18'b000000100100010100;
    n19324[771] = 18'b000000011100001100;
    n19324[770] = 18'b000000010100000110;
    n19324[769] = 18'b000000001100000010;
    n19324[768] = 18'b000000000100000000;
    n19324[767] = 18'b111111111000000000;
    n19324[766] = 18'b111111101000000110;
    n19324[765] = 18'b111111011000010010;
    n19324[764] = 18'b111111001000100100;
    n19324[763] = 18'b111110111000111010;
    n19324[762] = 18'b111110101001011000;
    n19324[761] = 18'b111110011001111100;
    n19324[760] = 18'b111110001010100100;
    n19324[759] = 18'b111101111011010010;
    n19324[758] = 18'b111101101100000110;
    n19324[757] = 18'b111101011100111110;
    n19324[756] = 18'b111101001101111110;
    n19324[755] = 18'b111100111111000010;
    n19324[754] = 18'b111100110000001010;
    n19324[753] = 18'b111100100001011010;
    n19324[752] = 18'b111100010010101110;
    n19324[751] = 18'b111100000100000110;
    n19324[750] = 18'b111011110101100100;
    n19324[749] = 18'b111011100111001000;
    n19324[748] = 18'b111011011000110000;
    n19324[747] = 18'b111011001010011110;
    n19324[746] = 18'b111010111100010000;
    n19324[745] = 18'b111010101110000110;
    n19324[744] = 18'b111010100000000010;
    n19324[743] = 18'b111010010010000100;
    n19324[742] = 18'b111010000100001000;
    n19324[741] = 18'b111001110110010100;
    n19324[740] = 18'b111001101000100010;
    n19324[739] = 18'b111001011010110110;
    n19324[738] = 18'b111001001101001110;
    n19324[737] = 18'b111000111111101010;
    n19324[736] = 18'b111000110010001100;
    n19324[735] = 18'b111000100100110010;
    n19324[734] = 18'b111000010111011100;
    n19324[733] = 18'b111000001010001010;
    n19324[732] = 18'b110111111100111110;
    n19324[731] = 18'b110111101111110110;
    n19324[730] = 18'b110111100010110010;
    n19324[729] = 18'b110111010101110010;
    n19324[728] = 18'b110111001000110110;
    n19324[727] = 18'b110110111011111110;
    n19324[726] = 18'b110110101111001010;
    n19324[725] = 18'b110110100010011010;
    n19324[724] = 18'b110110010101110000;
    n19324[723] = 18'b110110001001001000;
    n19324[722] = 18'b110101111100100110;
    n19324[721] = 18'b110101110000000110;
    n19324[720] = 18'b110101100011101010;
    n19324[719] = 18'b110101010111010100;
    n19324[718] = 18'b110101001011000000;
    n19324[717] = 18'b110100111110110000;
    n19324[716] = 18'b110100110010100100;
    n19324[715] = 18'b110100100110011100;
    n19324[714] = 18'b110100011010011000;
    n19324[713] = 18'b110100001110011000;
    n19324[712] = 18'b110100000010011100;
    n19324[711] = 18'b110011110110100010;
    n19324[710] = 18'b110011101010101100;
    n19324[709] = 18'b110011011110111100;
    n19324[708] = 18'b110011010011001100;
    n19324[707] = 18'b110011000111100010;
    n19324[706] = 18'b110010111011111100;
    n19324[705] = 18'b110010110000011000;
    n19324[704] = 18'b110010100100111000;
    n19324[703] = 18'b110010011001011010;
    n19324[702] = 18'b110010001110000010;
    n19324[701] = 18'b110010000010101100;
    n19324[700] = 18'b110001110111011000;
    n19324[699] = 18'b110001101100001010;
    n19324[698] = 18'b110001100000111110;
    n19324[697] = 18'b110001010101110110;
    n19324[696] = 18'b110001001010110000;
    n19324[695] = 18'b110000111111101110;
    n19324[694] = 18'b110000110100101110;
    n19324[693] = 18'b110000101001110100;
    n19324[692] = 18'b110000011110111010;
    n19324[691] = 18'b110000010100000110;
    n19324[690] = 18'b110000001001010100;
    n19324[689] = 18'b101111111110100100;
    n19324[688] = 18'b101111110011111000;
    n19324[687] = 18'b101111101001001110;
    n19324[686] = 18'b101111011110101000;
    n19324[685] = 18'b101111010100000110;
    n19324[684] = 18'b101111001001100110;
    n19324[683] = 18'b101110111111001010;
    n19324[682] = 18'b101110110100101110;
    n19324[681] = 18'b101110101010011000;
    n19324[680] = 18'b101110100000000100;
    n19324[679] = 18'b101110010101110010;
    n19324[678] = 18'b101110001011100100;
    n19324[677] = 18'b101110000001011000;
    n19324[676] = 18'b101101110111001110;
    n19324[675] = 18'b101101101101001000;
    n19324[674] = 18'b101101100011000110;
    n19324[673] = 18'b101101011001000110;
    n19324[672] = 18'b101101001111001000;
    n19324[671] = 18'b101101000101001100;
    n19324[670] = 18'b101100111011010100;
    n19324[669] = 18'b101100110001011110;
    n19324[668] = 18'b101100100111101010;
    n19324[667] = 18'b101100011101111010;
    n19324[666] = 18'b101100010100001100;
    n19324[665] = 18'b101100001010100010;
    n19324[664] = 18'b101100000000111000;
    n19324[663] = 18'b101011110111010010;
    n19324[662] = 18'b101011101101110000;
    n19324[661] = 18'b101011100100001110;
    n19324[660] = 18'b101011011010110000;
    n19324[659] = 18'b101011010001010100;
    n19324[658] = 18'b101011000111111010;
    n19324[657] = 18'b101010111110100100;
    n19324[656] = 18'b101010110101001110;
    n19324[655] = 18'b101010101011111100;
    n19324[654] = 18'b101010100010101100;
    n19324[653] = 18'b101010011001100000;
    n19324[652] = 18'b101010010000010100;
    n19324[651] = 18'b101010000111001100;
    n19324[650] = 18'b101001111110000110;
    n19324[649] = 18'b101001110101000010;
    n19324[648] = 18'b101001101100000000;
    n19324[647] = 18'b101001100011000010;
    n19324[646] = 18'b101001011010000100;
    n19324[645] = 18'b101001010001001010;
    n19324[644] = 18'b101001001000010000;
    n19324[643] = 18'b101000111111011010;
    n19324[642] = 18'b101000110110100110;
    n19324[641] = 18'b101000101101110100;
    n19324[640] = 18'b101000100101000110;
    n19324[639] = 18'b101000011100011000;
    n19324[638] = 18'b101000010011101100;
    n19324[637] = 18'b101000001011000100;
    n19324[636] = 18'b101000000010011100;
    n19324[635] = 18'b100111111001111000;
    n19324[634] = 18'b100111110001010110;
    n19324[633] = 18'b100111101000110100;
    n19324[632] = 18'b100111100000010110;
    n19324[631] = 18'b100111010111111010;
    n19324[630] = 18'b100111001111100000;
    n19324[629] = 18'b100111000111001000;
    n19324[628] = 18'b100110111110110000;
    n19324[627] = 18'b100110110110011100;
    n19324[626] = 18'b100110101110001010;
    n19324[625] = 18'b100110100101111010;
    n19324[624] = 18'b100110011101101100;
    n19324[623] = 18'b100110010101100000;
    n19324[622] = 18'b100110001101010110;
    n19324[621] = 18'b100110000101001100;
    n19324[620] = 18'b100101111101000110;
    n19324[619] = 18'b100101110101000010;
    n19324[618] = 18'b100101101101000000;
    n19324[617] = 18'b100101100100111110;
    n19324[616] = 18'b100101011101000000;
    n19324[615] = 18'b100101010101000010;
    n19324[614] = 18'b100101001101001000;
    n19324[613] = 18'b100101000101001110;
    n19324[612] = 18'b100100111101011000;
    n19324[611] = 18'b100100110101100010;
    n19324[610] = 18'b100100101101101110;
    n19324[609] = 18'b100100100101111100;
    n19324[608] = 18'b100100011110001100;
    n19324[607] = 18'b100100010110011110;
    n19324[606] = 18'b100100001110110000;
    n19324[605] = 18'b100100000111000110;
    n19324[604] = 18'b100011111111011110;
    n19324[603] = 18'b100011110111110110;
    n19324[602] = 18'b100011110000010000;
    n19324[601] = 18'b100011101000101100;
    n19324[600] = 18'b100011100001001010;
    n19324[599] = 18'b100011011001101010;
    n19324[598] = 18'b100011010010001100;
    n19324[597] = 18'b100011001010101110;
    n19324[596] = 18'b100011000011010010;
    n19324[595] = 18'b100010111011111010;
    n19324[594] = 18'b100010110100100000;
    n19324[593] = 18'b100010101101001010;
    n19324[592] = 18'b100010100101110110;
    n19324[591] = 18'b100010011110100010;
    n19324[590] = 18'b100010010111010010;
    n19324[589] = 18'b100010010000000010;
    n19324[588] = 18'b100010001000110100;
    n19324[587] = 18'b100010000001100110;
    n19324[586] = 18'b100001111010011100;
    n19324[585] = 18'b100001110011010010;
    n19324[584] = 18'b100001101100001010;
    n19324[583] = 18'b100001100101000100;
    n19324[582] = 18'b100001011101111110;
    n19324[581] = 18'b100001010110111010;
    n19324[580] = 18'b100001001111111010;
    n19324[579] = 18'b100001001000111000;
    n19324[578] = 18'b100001000001111010;
    n19324[577] = 18'b100000111010111100;
    n19324[576] = 18'b100000110100000000;
    n19324[575] = 18'b100000101101000110;
    n19324[574] = 18'b100000100110001110;
    n19324[573] = 18'b100000011111010110;
    n19324[572] = 18'b100000011000100000;
    n19324[571] = 18'b100000010001101100;
    n19324[570] = 18'b100000001010111000;
    n19324[569] = 18'b100000000100001000;
    n19324[568] = 18'b011111111101011000;
    n19324[567] = 18'b011111110110101000;
    n19324[566] = 18'b011111101111111100;
    n19324[565] = 18'b011111101001010000;
    n19324[564] = 18'b011111100010100100;
    n19324[563] = 18'b011111011011111100;
    n19324[562] = 18'b011111010101010100;
    n19324[561] = 18'b011111001110101110;
    n19324[560] = 18'b011111001000001000;
    n19324[559] = 18'b011111000001100100;
    n19324[558] = 18'b011110111011000010;
    n19324[557] = 18'b011110110100100010;
    n19324[556] = 18'b011110101110000010;
    n19324[555] = 18'b011110100111100100;
    n19324[554] = 18'b011110100001000110;
    n19324[553] = 18'b011110011010101010;
    n19324[552] = 18'b011110010100010000;
    n19324[551] = 18'b011110001101111000;
    n19324[550] = 18'b011110000111100000;
    n19324[549] = 18'b011110000001001010;
    n19324[548] = 18'b011101111010110100;
    n19324[547] = 18'b011101110100100000;
    n19324[546] = 18'b011101101110001110;
    n19324[545] = 18'b011101100111111100;
    n19324[544] = 18'b011101100001101100;
    n19324[543] = 18'b011101011011011110;
    n19324[542] = 18'b011101010101010000;
    n19324[541] = 18'b011101001111000100;
    n19324[540] = 18'b011101001000111000;
    n19324[539] = 18'b011101000010101110;
    n19324[538] = 18'b011100111100100110;
    n19324[537] = 18'b011100110110011110;
    n19324[536] = 18'b011100110000011000;
    n19324[535] = 18'b011100101010010100;
    n19324[534] = 18'b011100100100010000;
    n19324[533] = 18'b011100011110001100;
    n19324[532] = 18'b011100011000001010;
    n19324[531] = 18'b011100010010001010;
    n19324[530] = 18'b011100001100001100;
    n19324[529] = 18'b011100000110001110;
    n19324[528] = 18'b011100000000010000;
    n19324[527] = 18'b011011111010010100;
    n19324[526] = 18'b011011110100011010;
    n19324[525] = 18'b011011101110100000;
    n19324[524] = 18'b011011101000101000;
    n19324[523] = 18'b011011100010110010;
    n19324[522] = 18'b011011011100111100;
    n19324[521] = 18'b011011010111000110;
    n19324[520] = 18'b011011010001010010;
    n19324[519] = 18'b011011001011100000;
    n19324[518] = 18'b011011000101101110;
    n19324[517] = 18'b011010111111111110;
    n19324[516] = 18'b011010111010001110;
    n19324[515] = 18'b011010110100100000;
    n19324[514] = 18'b011010101110110100;
    n19324[513] = 18'b011010101001000110;
    n19324[512] = 18'b011010100011011100;
    n19324[511] = 18'b011010011101110010;
    n19324[510] = 18'b011010011000001000;
    n19324[509] = 18'b011010010010100000;
    n19324[508] = 18'b011010001100111010;
    n19324[507] = 18'b011010000111010100;
    n19324[506] = 18'b011010000001110000;
    n19324[505] = 18'b011001111100001100;
    n19324[504] = 18'b011001110110101000;
    n19324[503] = 18'b011001110001001000;
    n19324[502] = 18'b011001101011100110;
    n19324[501] = 18'b011001100110000110;
    n19324[500] = 18'b011001100000101000;
    n19324[499] = 18'b011001011011001010;
    n19324[498] = 18'b011001010101101110;
    n19324[497] = 18'b011001010000010010;
    n19324[496] = 18'b011001001010111000;
    n19324[495] = 18'b011001000101011110;
    n19324[494] = 18'b011001000000000100;
    n19324[493] = 18'b011000111010101110;
    n19324[492] = 18'b011000110101010110;
    n19324[491] = 18'b011000110000000000;
    n19324[490] = 18'b011000101010101100;
    n19324[489] = 18'b011000100101011000;
    n19324[488] = 18'b011000100000000100;
    n19324[487] = 18'b011000011010110010;
    n19324[486] = 18'b011000010101100010;
    n19324[485] = 18'b011000010000010010;
    n19324[484] = 18'b011000001011000010;
    n19324[483] = 18'b011000000101110100;
    n19324[482] = 18'b011000000000100110;
    n19324[481] = 18'b010111111011011010;
    n19324[480] = 18'b010111110110001110;
    n19324[479] = 18'b010111110001000100;
    n19324[478] = 18'b010111101011111010;
    n19324[477] = 18'b010111100110110010;
    n19324[476] = 18'b010111100001101010;
    n19324[475] = 18'b010111011100100100;
    n19324[474] = 18'b010111010111011110;
    n19324[473] = 18'b010111010010011000;
    n19324[472] = 18'b010111001101010100;
    n19324[471] = 18'b010111001000010000;
    n19324[470] = 18'b010111000011001110;
    n19324[469] = 18'b010110111110001100;
    n19324[468] = 18'b010110111001001100;
    n19324[467] = 18'b010110110100001100;
    n19324[466] = 18'b010110101111001100;
    n19324[465] = 18'b010110101010001110;
    n19324[464] = 18'b010110100101010000;
    n19324[463] = 18'b010110100000010100;
    n19324[462] = 18'b010110011011011000;
    n19324[461] = 18'b010110010110011110;
    n19324[460] = 18'b010110010001100100;
    n19324[459] = 18'b010110001100101010;
    n19324[458] = 18'b010110000111110010;
    n19324[457] = 18'b010110000010111010;
    n19324[456] = 18'b010101111110000100;
    n19324[455] = 18'b010101111001001110;
    n19324[454] = 18'b010101110100011010;
    n19324[453] = 18'b010101101111100110;
    n19324[452] = 18'b010101101010110010;
    n19324[451] = 18'b010101100110000000;
    n19324[450] = 18'b010101100001001110;
    n19324[449] = 18'b010101011100011100;
    n19324[448] = 18'b010101010111101100;
    n19324[447] = 18'b010101010010111100;
    n19324[446] = 18'b010101001110001110;
    n19324[445] = 18'b010101001001100000;
    n19324[444] = 18'b010101000100110100;
    n19324[443] = 18'b010101000000000110;
    n19324[442] = 18'b010100111011011100;
    n19324[441] = 18'b010100110110110000;
    n19324[440] = 18'b010100110010000110;
    n19324[439] = 18'b010100101101011110;
    n19324[438] = 18'b010100101000110110;
    n19324[437] = 18'b010100100100001110;
    n19324[436] = 18'b010100011111100110;
    n19324[435] = 18'b010100011011000000;
    n19324[434] = 18'b010100010110011010;
    n19324[433] = 18'b010100010001110110;
    n19324[432] = 18'b010100001101010010;
    n19324[431] = 18'b010100001000110000;
    n19324[430] = 18'b010100000100001100;
    n19324[429] = 18'b010011111111101010;
    n19324[428] = 18'b010011111011001010;
    n19324[427] = 18'b010011110110101010;
    n19324[426] = 18'b010011110010001010;
    n19324[425] = 18'b010011101101101100;
    n19324[424] = 18'b010011101001001110;
    n19324[423] = 18'b010011100100110000;
    n19324[422] = 18'b010011100000010100;
    n19324[421] = 18'b010011011011111000;
    n19324[420] = 18'b010011010111011100;
    n19324[419] = 18'b010011010011000010;
    n19324[418] = 18'b010011001110101000;
    n19324[417] = 18'b010011001010001110;
    n19324[416] = 18'b010011000101110110;
    n19324[415] = 18'b010011000001011110;
    n19324[414] = 18'b010010111101001000;
    n19324[413] = 18'b010010111000110000;
    n19324[412] = 18'b010010110100011010;
    n19324[411] = 18'b010010110000000110;
    n19324[410] = 18'b010010101011110010;
    n19324[409] = 18'b010010100111011110;
    n19324[408] = 18'b010010100011001010;
    n19324[407] = 18'b010010011110111000;
    n19324[406] = 18'b010010011010100110;
    n19324[405] = 18'b010010010110010110;
    n19324[404] = 18'b010010010010000110;
    n19324[403] = 18'b010010001101110110;
    n19324[402] = 18'b010010001001100110;
    n19324[401] = 18'b010010000101011000;
    n19324[400] = 18'b010010000001001010;
    n19324[399] = 18'b010001111100111110;
    n19324[398] = 18'b010001111000110010;
    n19324[397] = 18'b010001110100100110;
    n19324[396] = 18'b010001110000011010;
    n19324[395] = 18'b010001101100010000;
    n19324[394] = 18'b010001101000000110;
    n19324[393] = 18'b010001100011111100;
    n19324[392] = 18'b010001011111110100;
    n19324[391] = 18'b010001011011101100;
    n19324[390] = 18'b010001010111100100;
    n19324[389] = 18'b010001010011011110;
    n19324[388] = 18'b010001001111011000;
    n19324[387] = 18'b010001001011010010;
    n19324[386] = 18'b010001000111001110;
    n19324[385] = 18'b010001000011001010;
    n19324[384] = 18'b010000111111000110;
    n19324[383] = 18'b010000111011000010;
    n19324[382] = 18'b010000110111000000;
    n19324[381] = 18'b010000110010111110;
    n19324[380] = 18'b010000101110111100;
    n19324[379] = 18'b010000101010111100;
    n19324[378] = 18'b010000100110111100;
    n19324[377] = 18'b010000100010111100;
    n19324[376] = 18'b010000011110111110;
    n19324[375] = 18'b010000011011000000;
    n19324[374] = 18'b010000010111000010;
    n19324[373] = 18'b010000010011000100;
    n19324[372] = 18'b010000001111001000;
    n19324[371] = 18'b010000001011001100;
    n19324[370] = 18'b010000000111010000;
    n19324[369] = 18'b010000000011010110;
    n19324[368] = 18'b001111111111011100;
    n19324[367] = 18'b001111111011100010;
    n19324[366] = 18'b001111110111101010;
    n19324[365] = 18'b001111110011110000;
    n19324[364] = 18'b001111101111111000;
    n19324[363] = 18'b001111101100000010;
    n19324[362] = 18'b001111101000001010;
    n19324[361] = 18'b001111100100010100;
    n19324[360] = 18'b001111100000011110;
    n19324[359] = 18'b001111011100101010;
    n19324[358] = 18'b001111011000110110;
    n19324[357] = 18'b001111010101000010;
    n19324[356] = 18'b001111010001001110;
    n19324[355] = 18'b001111001101011010;
    n19324[354] = 18'b001111001001101000;
    n19324[353] = 18'b001111000101110110;
    n19324[352] = 18'b001111000010000110;
    n19324[351] = 18'b001110111110010100;
    n19324[350] = 18'b001110111010100100;
    n19324[349] = 18'b001110110110110100;
    n19324[348] = 18'b001110110011000110;
    n19324[347] = 18'b001110101111010110;
    n19324[346] = 18'b001110101011101000;
    n19324[345] = 18'b001110100111111010;
    n19324[344] = 18'b001110100100001110;
    n19324[343] = 18'b001110100000100010;
    n19324[342] = 18'b001110011100110110;
    n19324[341] = 18'b001110011001001010;
    n19324[340] = 18'b001110010101011110;
    n19324[339] = 18'b001110010001110100;
    n19324[338] = 18'b001110001110001010;
    n19324[337] = 18'b001110001010100000;
    n19324[336] = 18'b001110000110111000;
    n19324[335] = 18'b001110000011010000;
    n19324[334] = 18'b001101111111101000;
    n19324[333] = 18'b001101111100000000;
    n19324[332] = 18'b001101111000011010;
    n19324[331] = 18'b001101110100110010;
    n19324[330] = 18'b001101110001001100;
    n19324[329] = 18'b001101101101101000;
    n19324[328] = 18'b001101101010000010;
    n19324[327] = 18'b001101100110011110;
    n19324[326] = 18'b001101100010111010;
    n19324[325] = 18'b001101011111010110;
    n19324[324] = 18'b001101011011110100;
    n19324[323] = 18'b001101011000010010;
    n19324[322] = 18'b001101010100110000;
    n19324[321] = 18'b001101010001001110;
    n19324[320] = 18'b001101001101101100;
    n19324[319] = 18'b001101001010001100;
    n19324[318] = 18'b001101000110101100;
    n19324[317] = 18'b001101000011001100;
    n19324[316] = 18'b001100111111101110;
    n19324[315] = 18'b001100111100001110;
    n19324[314] = 18'b001100111000110000;
    n19324[313] = 18'b001100110101010100;
    n19324[312] = 18'b001100110001110110;
    n19324[311] = 18'b001100101110011010;
    n19324[310] = 18'b001100101010111100;
    n19324[309] = 18'b001100100111100000;
    n19324[308] = 18'b001100100100000110;
    n19324[307] = 18'b001100100000101010;
    n19324[306] = 18'b001100011101010000;
    n19324[305] = 18'b001100011001110110;
    n19324[304] = 18'b001100010110011100;
    n19324[303] = 18'b001100010011000100;
    n19324[302] = 18'b001100001111101010;
    n19324[301] = 18'b001100001100010010;
    n19324[300] = 18'b001100001000111010;
    n19324[299] = 18'b001100000101100100;
    n19324[298] = 18'b001100000010001100;
    n19324[297] = 18'b001011111110110110;
    n19324[296] = 18'b001011111011100000;
    n19324[295] = 18'b001011111000001010;
    n19324[294] = 18'b001011110100110110;
    n19324[293] = 18'b001011110001100010;
    n19324[292] = 18'b001011101110001100;
    n19324[291] = 18'b001011101010111010;
    n19324[290] = 18'b001011100111100110;
    n19324[289] = 18'b001011100100010010;
    n19324[288] = 18'b001011100001000000;
    n19324[287] = 18'b001011011101101110;
    n19324[286] = 18'b001011011010011100;
    n19324[285] = 18'b001011010111001100;
    n19324[284] = 18'b001011010011111010;
    n19324[283] = 18'b001011010000101010;
    n19324[282] = 18'b001011001101011010;
    n19324[281] = 18'b001011001010001010;
    n19324[280] = 18'b001011000110111100;
    n19324[279] = 18'b001011000011101110;
    n19324[278] = 18'b001011000000011110;
    n19324[277] = 18'b001010111101010000;
    n19324[276] = 18'b001010111010000100;
    n19324[275] = 18'b001010110110110110;
    n19324[274] = 18'b001010110011101010;
    n19324[273] = 18'b001010110000011110;
    n19324[272] = 18'b001010101101010010;
    n19324[271] = 18'b001010101010000110;
    n19324[270] = 18'b001010100110111100;
    n19324[269] = 18'b001010100011110000;
    n19324[268] = 18'b001010100000100110;
    n19324[267] = 18'b001010011101011100;
    n19324[266] = 18'b001010011010010100;
    n19324[265] = 18'b001010010111001010;
    n19324[264] = 18'b001010010100000010;
    n19324[263] = 18'b001010010000111010;
    n19324[262] = 18'b001010001101110010;
    n19324[261] = 18'b001010001010101010;
    n19324[260] = 18'b001010000111100100;
    n19324[259] = 18'b001010000100011100;
    n19324[258] = 18'b001010000001010110;
    n19324[257] = 18'b001001111110010000;
    n19324[256] = 18'b001001111011001100;
    n19324[255] = 18'b001001111000000110;
    n19324[254] = 18'b001001110101000010;
    n19324[253] = 18'b001001110001111110;
    n19324[252] = 18'b001001101110111010;
    n19324[251] = 18'b001001101011110110;
    n19324[250] = 18'b001001101000110010;
    n19324[249] = 18'b001001100101110000;
    n19324[248] = 18'b001001100010101110;
    n19324[247] = 18'b001001011111101100;
    n19324[246] = 18'b001001011100101010;
    n19324[245] = 18'b001001011001101000;
    n19324[244] = 18'b001001010110101000;
    n19324[243] = 18'b001001010011101000;
    n19324[242] = 18'b001001010000100110;
    n19324[241] = 18'b001001001101101000;
    n19324[240] = 18'b001001001010101000;
    n19324[239] = 18'b001001000111101000;
    n19324[238] = 18'b001001000100101010;
    n19324[237] = 18'b001001000001101100;
    n19324[236] = 18'b001000111110101110;
    n19324[235] = 18'b001000111011110000;
    n19324[234] = 18'b001000111000110010;
    n19324[233] = 18'b001000110101110110;
    n19324[232] = 18'b001000110010111010;
    n19324[231] = 18'b001000101111111110;
    n19324[230] = 18'b001000101101000010;
    n19324[229] = 18'b001000101010000110;
    n19324[228] = 18'b001000100111001010;
    n19324[227] = 18'b001000100100010000;
    n19324[226] = 18'b001000100001010110;
    n19324[225] = 18'b001000011110011100;
    n19324[224] = 18'b001000011011100010;
    n19324[223] = 18'b001000011000101000;
    n19324[222] = 18'b001000010101110000;
    n19324[221] = 18'b001000010010110110;
    n19324[220] = 18'b001000001111111110;
    n19324[219] = 18'b001000001101000110;
    n19324[218] = 18'b001000001010001110;
    n19324[217] = 18'b001000000111011000;
    n19324[216] = 18'b001000000100100000;
    n19324[215] = 18'b001000000001101010;
    n19324[214] = 18'b000111111110110100;
    n19324[213] = 18'b000111111011111110;
    n19324[212] = 18'b000111111001001000;
    n19324[211] = 18'b000111110110010010;
    n19324[210] = 18'b000111110011011110;
    n19324[209] = 18'b000111110000101010;
    n19324[208] = 18'b000111101101110110;
    n19324[207] = 18'b000111101011000010;
    n19324[206] = 18'b000111101000001110;
    n19324[205] = 18'b000111100101011010;
    n19324[204] = 18'b000111100010101000;
    n19324[203] = 18'b000111011111110100;
    n19324[202] = 18'b000111011101000010;
    n19324[201] = 18'b000111011010010000;
    n19324[200] = 18'b000111010111011110;
    n19324[199] = 18'b000111010100101110;
    n19324[198] = 18'b000111010001111100;
    n19324[197] = 18'b000111001111001100;
    n19324[196] = 18'b000111001100011100;
    n19324[195] = 18'b000111001001101100;
    n19324[194] = 18'b000111000110111100;
    n19324[193] = 18'b000111000100001100;
    n19324[192] = 18'b000111000001011110;
    n19324[191] = 18'b000110111110101110;
    n19324[190] = 18'b000110111100000000;
    n19324[189] = 18'b000110111001010010;
    n19324[188] = 18'b000110110110100100;
    n19324[187] = 18'b000110110011110110;
    n19324[186] = 18'b000110110001001010;
    n19324[185] = 18'b000110101110011100;
    n19324[184] = 18'b000110101011110000;
    n19324[183] = 18'b000110101001000100;
    n19324[182] = 18'b000110100110011000;
    n19324[181] = 18'b000110100011101100;
    n19324[180] = 18'b000110100001000000;
    n19324[179] = 18'b000110011110010110;
    n19324[178] = 18'b000110011011101010;
    n19324[177] = 18'b000110011001000000;
    n19324[176] = 18'b000110010110010110;
    n19324[175] = 18'b000110010011101100;
    n19324[174] = 18'b000110010001000010;
    n19324[173] = 18'b000110001110011010;
    n19324[172] = 18'b000110001011110000;
    n19324[171] = 18'b000110001001001000;
    n19324[170] = 18'b000110000110100000;
    n19324[169] = 18'b000110000011111000;
    n19324[168] = 18'b000110000001010000;
    n19324[167] = 18'b000101111110101000;
    n19324[166] = 18'b000101111100000000;
    n19324[165] = 18'b000101111001011010;
    n19324[164] = 18'b000101110110110100;
    n19324[163] = 18'b000101110100001110;
    n19324[162] = 18'b000101110001101000;
    n19324[161] = 18'b000101101111000010;
    n19324[160] = 18'b000101101100011100;
    n19324[159] = 18'b000101101001110110;
    n19324[158] = 18'b000101100111010010;
    n19324[157] = 18'b000101100100101110;
    n19324[156] = 18'b000101100010001000;
    n19324[155] = 18'b000101011111100100;
    n19324[154] = 18'b000101011101000010;
    n19324[153] = 18'b000101011010011110;
    n19324[152] = 18'b000101010111111010;
    n19324[151] = 18'b000101010101011000;
    n19324[150] = 18'b000101010010110110;
    n19324[149] = 18'b000101010000010010;
    n19324[148] = 18'b000101001101110000;
    n19324[147] = 18'b000101001011001110;
    n19324[146] = 18'b000101001000101110;
    n19324[145] = 18'b000101000110001100;
    n19324[144] = 18'b000101000011101100;
    n19324[143] = 18'b000101000001001010;
    n19324[142] = 18'b000100111110101010;
    n19324[141] = 18'b000100111100001010;
    n19324[140] = 18'b000100111001101010;
    n19324[139] = 18'b000100110111001010;
    n19324[138] = 18'b000100110100101100;
    n19324[137] = 18'b000100110010001100;
    n19324[136] = 18'b000100101111101110;
    n19324[135] = 18'b000100101101010000;
    n19324[134] = 18'b000100101010110000;
    n19324[133] = 18'b000100101000010010;
    n19324[132] = 18'b000100100101110110;
    n19324[131] = 18'b000100100011011000;
    n19324[130] = 18'b000100100000111010;
    n19324[129] = 18'b000100011110011110;
    n19324[128] = 18'b000100011100000000;
    n19324[127] = 18'b000100011001100100;
    n19324[126] = 18'b000100010111001000;
    n19324[125] = 18'b000100010100101100;
    n19324[124] = 18'b000100010010010000;
    n19324[123] = 18'b000100001111110110;
    n19324[122] = 18'b000100001101011010;
    n19324[121] = 18'b000100001011000000;
    n19324[120] = 18'b000100001000100110;
    n19324[119] = 18'b000100000110001010;
    n19324[118] = 18'b000100000011110000;
    n19324[117] = 18'b000100000001010110;
    n19324[116] = 18'b000011111110111110;
    n19324[115] = 18'b000011111100100100;
    n19324[114] = 18'b000011111010001100;
    n19324[113] = 18'b000011110111110010;
    n19324[112] = 18'b000011110101011010;
    n19324[111] = 18'b000011110011000010;
    n19324[110] = 18'b000011110000101010;
    n19324[109] = 18'b000011101110010010;
    n19324[108] = 18'b000011101011111010;
    n19324[107] = 18'b000011101001100010;
    n19324[106] = 18'b000011100111001100;
    n19324[105] = 18'b000011100100110100;
    n19324[104] = 18'b000011100010011110;
    n19324[103] = 18'b000011100000001000;
    n19324[102] = 18'b000011011101110010;
    n19324[101] = 18'b000011011011011100;
    n19324[100] = 18'b000011011001000110;
    n19324[99] = 18'b000011010110110010;
    n19324[98] = 18'b000011010100011100;
    n19324[97] = 18'b000011010010001000;
    n19324[96] = 18'b000011001111110010;
    n19324[95] = 18'b000011001101011110;
    n19324[94] = 18'b000011001011001010;
    n19324[93] = 18'b000011001000110110;
    n19324[92] = 18'b000011000110100010;
    n19324[91] = 18'b000011000100010000;
    n19324[90] = 18'b000011000001111100;
    n19324[89] = 18'b000010111111101010;
    n19324[88] = 18'b000010111101010110;
    n19324[87] = 18'b000010111011000100;
    n19324[86] = 18'b000010111000110010;
    n19324[85] = 18'b000010110110100000;
    n19324[84] = 18'b000010110100001110;
    n19324[83] = 18'b000010110001111100;
    n19324[82] = 18'b000010101111101100;
    n19324[81] = 18'b000010101101011010;
    n19324[80] = 18'b000010101011001010;
    n19324[79] = 18'b000010101000111000;
    n19324[78] = 18'b000010100110101000;
    n19324[77] = 18'b000010100100011000;
    n19324[76] = 18'b000010100010001000;
    n19324[75] = 18'b000010011111111000;
    n19324[74] = 18'b000010011101101010;
    n19324[73] = 18'b000010011011011010;
    n19324[72] = 18'b000010011001001010;
    n19324[71] = 18'b000010010110111100;
    n19324[70] = 18'b000010010100101110;
    n19324[69] = 18'b000010010010100000;
    n19324[68] = 18'b000010010000010000;
    n19324[67] = 18'b000010001110000100;
    n19324[66] = 18'b000010001011110110;
    n19324[65] = 18'b000010001001101000;
    n19324[64] = 18'b000010000111011010;
    n19324[63] = 18'b000010000101001110;
    n19324[62] = 18'b000010000011000000;
    n19324[61] = 18'b000010000000110100;
    n19324[60] = 18'b000001111110101000;
    n19324[59] = 18'b000001111100011100;
    n19324[58] = 18'b000001111010010000;
    n19324[57] = 18'b000001111000000100;
    n19324[56] = 18'b000001110101111000;
    n19324[55] = 18'b000001110011101110;
    n19324[54] = 18'b000001110001100010;
    n19324[53] = 18'b000001101111011000;
    n19324[52] = 18'b000001101101001100;
    n19324[51] = 18'b000001101011000010;
    n19324[50] = 18'b000001101000111000;
    n19324[49] = 18'b000001100110101110;
    n19324[48] = 18'b000001100100100100;
    n19324[47] = 18'b000001100010011100;
    n19324[46] = 18'b000001100000010010;
    n19324[45] = 18'b000001011110001000;
    n19324[44] = 18'b000001011100000000;
    n19324[43] = 18'b000001011001110110;
    n19324[42] = 18'b000001010111101110;
    n19324[41] = 18'b000001010101100110;
    n19324[40] = 18'b000001010011011110;
    n19324[39] = 18'b000001010001010110;
    n19324[38] = 18'b000001001111001110;
    n19324[37] = 18'b000001001101000110;
    n19324[36] = 18'b000001001011000000;
    n19324[35] = 18'b000001001000111000;
    n19324[34] = 18'b000001000110110010;
    n19324[33] = 18'b000001000100101100;
    n19324[32] = 18'b000001000010100100;
    n19324[31] = 18'b000001000000011110;
    n19324[30] = 18'b000000111110011000;
    n19324[29] = 18'b000000111100010010;
    n19324[28] = 18'b000000111010001100;
    n19324[27] = 18'b000000111000001000;
    n19324[26] = 18'b000000110110000010;
    n19324[25] = 18'b000000110011111110;
    n19324[24] = 18'b000000110001111000;
    n19324[23] = 18'b000000101111110100;
    n19324[22] = 18'b000000101101110000;
    n19324[21] = 18'b000000101011101100;
    n19324[20] = 18'b000000101001101000;
    n19324[19] = 18'b000000100111100100;
    n19324[18] = 18'b000000100101100000;
    n19324[17] = 18'b000000100011011100;
    n19324[16] = 18'b000000100001011000;
    n19324[15] = 18'b000000011111010110;
    n19324[14] = 18'b000000011101010010;
    n19324[13] = 18'b000000011011010000;
    n19324[12] = 18'b000000011001001110;
    n19324[11] = 18'b000000010111001100;
    n19324[10] = 18'b000000010101001010;
    n19324[9] = 18'b000000010011001000;
    n19324[8] = 18'b000000010001000110;
    n19324[7] = 18'b000000001111000100;
    n19324[6] = 18'b000000001101000010;
    n19324[5] = 18'b000000001011000010;
    n19324[4] = 18'b000000001001000000;
    n19324[3] = 18'b000000000111000000;
    n19324[2] = 18'b000000000101000000;
    n19324[1] = 18'b000000000011000000;
    n19324[0] = 18'b000000000001000000;
    end
  assign n19325_data = n19324[n13032_o];
  /* fpu.vhdl:571:48  */
endmodule

module execute1_0_47ec8d98366433dc002e7721c9e37d5067547937
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  clk,
   input  rst,
   input  flush_in,
   input  e_in_valid,
   input  [1:0] e_in_unit,
   input  e_in_fac,
   input  [5:0] e_in_insn_type,
   input  [63:0] e_in_nia,
   input  [2:0] e_in_instr_tag,
   input  [6:0] e_in_write_reg,
   input  e_in_write_reg_enable,
   input  [6:0] e_in_read_reg1,
   input  [6:0] e_in_read_reg2,
   input  [63:0] e_in_read_data1,
   input  [63:0] e_in_read_data2,
   input  [63:0] e_in_read_data3,
   input  [31:0] e_in_cr,
   input  [4:0] e_in_xerc,
   input  e_in_lr,
   input  e_in_br_abs,
   input  e_in_rc,
   input  e_in_oe,
   input  e_in_invert_a,
   input  e_in_addm1,
   input  e_in_invert_out,
   input  [1:0] e_in_input_carry,
   input  e_in_output_carry,
   input  e_in_input_cr,
   input  e_in_output_cr,
   input  e_in_output_xer,
   input  e_in_is_32bit,
   input  e_in_is_signed,
   input  [31:0] e_in_insn,
   input  [3:0] e_in_data_len,
   input  e_in_byte_reverse,
   input  e_in_sign_extend,
   input  e_in_update,
   input  e_in_reserve,
   input  e_in_br_pred,
   input  [2:0] e_in_result_sel,
   input  [2:0] e_in_sub_select,
   input  e_in_repeat,
   input  e_in_second,
   input  l_in_busy,
   input  l_in_in_progress,
   input  l_in_interrupt,
   input  fp_in_busy,
   input  fp_in_exception,
   input  ext_irq_in,
   input  interrupt_in,
   input  wb_events_instr_complete,
   input  wb_events_fp_complete,
   input  ls_events_load_complete,
   input  ls_events_store_complete,
   input  ls_events_itlb_miss,
   input  dc_events_load_miss,
   input  dc_events_store_miss,
   input  dc_events_dcache_refill,
   input  dc_events_dtlb_miss,
   input  dc_events_dtlb_miss_resolved,
   input  ic_events_icache_miss,
   input  ic_events_itlb_miss_resolved,
   input  [63:0] log_rd_data,
   input  [31:0] log_wr_addr,
   output busy_out,
   output l_out_valid,
   output [5:0] l_out_op,
   output [63:0] l_out_nia,
   output [31:0] l_out_insn,
   output [2:0] l_out_instr_tag,
   output [63:0] l_out_addr1,
   output [63:0] l_out_addr2,
   output [63:0] l_out_data,
   output [6:0] l_out_write_reg,
   output [3:0] l_out_length,
   output l_out_ci,
   output l_out_byte_reverse,
   output l_out_sign_extend,
   output l_out_update,
   output [4:0] l_out_xerc,
   output l_out_reserve,
   output l_out_rc,
   output l_out_virt_mode,
   output l_out_priv_mode,
   output l_out_mode_32bit,
   output l_out_is_32bit,
   output l_out_repeat,
   output l_out_second,
   output [63:0] l_out_msr,
   output fp_out_valid,
   output [5:0] fp_out_op,
   output [63:0] fp_out_nia,
   output [2:0] fp_out_itag,
   output [31:0] fp_out_insn,
   output fp_out_single,
   output [1:0] fp_out_fe_mode,
   output [63:0] fp_out_fra,
   output [63:0] fp_out_frb,
   output [63:0] fp_out_frc,
   output [6:0] fp_out_frt,
   output fp_out_rc,
   output fp_out_out_cr,
   output e_out_valid,
   output [2:0] e_out_instr_tag,
   output e_out_rc,
   output e_out_mode_32bit,
   output e_out_write_enable,
   output [6:0] e_out_write_reg,
   output [63:0] e_out_write_data,
   output e_out_write_cr_enable,
   output [7:0] e_out_write_cr_mask,
   output [31:0] e_out_write_cr_data,
   output e_out_write_xerc_enable,
   output [4:0] e_out_xerc,
   output e_out_interrupt,
   output [11:0] e_out_intr_vec,
   output e_out_redirect,
   output [3:0] e_out_redir_mode,
   output [63:0] e_out_last_nia,
   output [63:0] e_out_br_offset,
   output e_out_br_last,
   output e_out_br_taken,
   output e_out_abs_br,
   output [15:0] e_out_srr1,
   output [63:0] e_out_msr,
   output [2:0] bypass_data_tag,
   output [63:0] bypass_data_data,
   output [2:0] bypass_cr_data_tag,
   output [31:0] bypass_cr_data_data,
   output [63:0] dbg_msr_out,
   output icache_inval,
   output terminate_out,
   output [14:0] log_out,
   output [31:0] log_rd_addr);
  wire [391:0] n9139_o;
  wire [2:0] n9140_o;
  wire [1:0] n9141_o;
  wire n9143_o;
  wire [5:0] n9144_o;
  wire [63:0] n9145_o;
  wire [31:0] n9146_o;
  wire [2:0] n9147_o;
  wire [63:0] n9148_o;
  wire [63:0] n9149_o;
  wire [63:0] n9150_o;
  wire [6:0] n9151_o;
  wire [3:0] n9152_o;
  wire n9153_o;
  wire n9154_o;
  wire n9155_o;
  wire n9156_o;
  wire [4:0] n9157_o;
  wire n9158_o;
  wire n9159_o;
  wire n9160_o;
  wire n9161_o;
  wire n9162_o;
  wire n9163_o;
  wire n9164_o;
  wire n9165_o;
  wire [63:0] n9166_o;
  wire n9168_o;
  wire [5:0] n9169_o;
  wire [63:0] n9170_o;
  wire [2:0] n9171_o;
  wire [31:0] n9172_o;
  wire n9173_o;
  wire [1:0] n9174_o;
  wire [63:0] n9175_o;
  wire [63:0] n9176_o;
  wire [63:0] n9177_o;
  wire [6:0] n9178_o;
  wire n9179_o;
  wire n9180_o;
  wire n9182_o;
  wire [2:0] n9183_o;
  wire n9184_o;
  wire n9185_o;
  wire n9186_o;
  wire [6:0] n9187_o;
  wire [63:0] n9188_o;
  wire n9189_o;
  wire [7:0] n9190_o;
  wire [31:0] n9191_o;
  wire n9192_o;
  wire [4:0] n9193_o;
  wire n9194_o;
  wire [11:0] n9195_o;
  wire n9196_o;
  wire [3:0] n9197_o;
  wire [63:0] n9198_o;
  wire [63:0] n9199_o;
  wire n9200_o;
  wire n9201_o;
  wire n9202_o;
  wire [15:0] n9203_o;
  wire [63:0] n9204_o;
  wire [2:0] n9206_o;
  wire [63:0] n9207_o;
  wire [2:0] n9209_o;
  wire [31:0] n9210_o;
  wire [1:0] n9214_o;
  wire [2:0] n9215_o;
  wire [4:0] n9216_o;
  wire [1:0] n9217_o;
  wire [798:0] r;
  wire [798:0] rin;
  wire [63:0] a_in;
  wire [63:0] b_in;
  wire [63:0] c_in;
  wire [31:0] cr_in;
  wire [4:0] xerc_in;
  wire valid_in;
  reg [255:0] ctrl;
  reg [255:0] ctrl_tmp;
  wire right_shift;
  wire rot_clear_left;
  wire rot_clear_right;
  wire rot_sign_ext;
  wire [63:0] rotator_result;
  wire rotator_carry;
  wire [63:0] logical_result;
  wire do_popcnt;
  wire [63:0] countbits_result;
  wire [63:0] alu_result;
  wire [63:0] adder_result;
  wire [63:0] misc_result;
  wire [63:0] muldiv_result;
  wire [63:0] spr_result;
  wire [63:0] next_nia;
  wire [391:0] current;
  wire carry_32;
  wire carry_64;
  wire overflow_32;
  wire overflow_64;
  wire [4:0] trapval;
  wire [7:0] write_cr_mask;
  wire [31:0] write_cr_data;
  wire [258:0] x_to_multiply;
  wire [129:0] multiply_to_x;
  wire [133:0] x_to_divider;
  wire [65:0] divider_to_x;
  wire [63:0] random_raw;
  wire [63:0] random_cond;
  wire random_err;
  wire [227:0] x_to_pmu;
  wire [64:0] pmu_to_x;
  wire [63:0] rotator_0_result;
  wire rotator_0_carry_out;
  wire [6:0] n9223_o;
  wire [31:0] n9224_o;
  wire n9225_o;
  wire n9226_o;
  wire [63:0] logical_0_result;
  wire [5:0] n9229_o;
  wire n9230_o;
  wire n9231_o;
  wire [3:0] n9233_o;
  wire [63:0] countbits_0_result;
  wire n9234_o;
  wire n9235_o;
  wire [3:0] n9236_o;
  wire multiply_0_m_out_valid;
  wire [127:0] multiply_0_m_out_result;
  wire multiply_0_m_out_overflow;
  wire n9238_o;
  wire [63:0] n9239_o;
  wire [63:0] n9240_o;
  wire [127:0] n9241_o;
  wire n9242_o;
  wire n9243_o;
  wire [129:0] n9244_o;
  wire divider_0_d_out_valid;
  wire [63:0] divider_0_d_out_write_reg_data;
  wire divider_0_d_out_overflow;
  wire n9246_o;
  wire [63:0] n9247_o;
  wire [63:0] n9248_o;
  wire n9249_o;
  wire n9250_o;
  wire n9251_o;
  wire n9252_o;
  wire n9253_o;
  wire [65:0] n9254_o;
  wire [63:0] random_0_data;
  wire [63:0] random_0_raw;
  wire random_0_err;
  wire [63:0] pmu_0_p_out_spr_val;
  wire pmu_0_p_out_intr;
  wire n9259_o;
  wire n9260_o;
  wire [4:0] n9261_o;
  wire [63:0] n9262_o;
  wire [3:0] n9263_o;
  wire n9264_o;
  wire n9265_o;
  wire n9266_o;
  wire [63:0] n9267_o;
  wire [63:0] n9268_o;
  wire n9269_o;
  wire [20:0] n9270_o;
  wire [64:0] n9271_o;
  wire [63:0] n9273_o;
  wire [31:0] n9274_o;
  wire [63:0] n9275_o;
  wire [63:0] n9276_o;
  wire [63:0] n9277_o;
  wire [31:0] n9278_o;
  wire n9279_o;
  wire n9280_o;
  wire n9281_o;
  wire n9282_o;
  wire n9283_o;
  wire n9284_o;
  wire n9285_o;
  wire n9286_o;
  wire n9287_o;
  wire n9288_o;
  wire n9289_o;
  wire n9290_o;
  wire n9291_o;
  wire n9292_o;
  wire n9293_o;
  wire n9294_o;
  wire n9295_o;
  wire [3:0] n9300_o;
  wire [3:0] n9301_o;
  wire [3:0] n9302_o;
  wire [3:0] n9303_o;
  wire [3:0] n9304_o;
  wire [15:0] n9305_o;
  wire [4:0] n9306_o;
  wire [20:0] n9307_o;
  wire [63:0] n9308_o;
  wire [4:0] n9311_o;
  wire [353:0] n9313_o;
  wire [4:0] n9314_o;
  wire [353:0] n9315_o;
  wire n9316_o;
  wire n9317_o;
  wire n9318_o;
  wire [4:0] n9319_o;
  wire [4:0] n9320_o;
  wire [1:0] n9321_o;
  wire n9322_o;
  wire n9323_o;
  wire n9324_o;
  wire n9325_o;
  wire n9326_o;
  wire n9328_o;
  wire n9329_o;
  wire n9330_o;
  wire n9331_o;
  wire n9332_o;
  wire n9333_o;
  wire n9334_o;
  wire n9335_o;
  reg n9336_o;
  wire n9337_o;
  wire n9338_o;
  wire n9339_o;
  wire n9340_o;
  wire n9341_o;
  wire n9342_o;
  wire n9343_o;
  wire n9344_o;
  wire [391:0] n9345_o;
  wire [391:0] n9346_o;
  wire [2:0] n9347_o;
  wire n9349_o;
  wire n9351_o;
  wire n9353_o;
  wire n9355_o;
  wire n9357_o;
  wire n9359_o;
  wire n9361_o;
  wire [6:0] n9362_o;
  reg [63:0] n9363_o;
  wire [798:0] n9370_o;
  wire [191:0] n9371_o;
  wire [191:0] n9372_o;
  wire [191:0] n9373_o;
  wire [63:0] n9374_o;
  wire [63:0] n9375_o;
  wire [63:0] n9376_o;
  wire [255:0] n9378_o;
  wire n9420_o;
  wire n9421_o;
  wire [63:0] n9422_o;
  wire [63:0] n9423_o;
  wire n9424_o;
  wire n9425_o;
  wire [63:0] n9427_o;
  wire [1:0] n9430_o;
  wire n9437_o;
  wire n9438_o;
  wire n9440_o;
  wire n9441_o;
  wire n9443_o;
  wire n9446_o;
  wire [3:0] n9447_o;
  reg n9449_o;
  wire [64:0] n9454_o;
  wire [64:0] n9455_o;
  wire [64:0] n9456_o;
  wire [64:0] n9457_o;
  wire [64:0] n9458_o;
  wire [63:0] n9459_o;
  wire n9460_o;
  wire n9461_o;
  wire n9462_o;
  wire n9463_o;
  wire n9464_o;
  wire n9465_o;
  wire n9467_o;
  wire n9468_o;
  wire n9469_o;
  wire n9474_o;
  wire n9475_o;
  wire n9476_o;
  wire n9477_o;
  wire n9479_o;
  wire n9480_o;
  wire n9481_o;
  wire n9486_o;
  wire n9487_o;
  wire n9488_o;
  wire n9489_o;
  wire n9490_o;
  wire n9491_o;
  wire n9492_o;
  wire n9493_o;
  wire n9494_o;
  wire n9495_o;
  wire n9496_o;
  wire n9497_o;
  wire n9499_o;
  wire n9502_o;
  wire n9504_o;
  wire [63:0] n9505_o;
  wire [63:0] n9506_o;
  wire n9507_o;
  wire [63:0] n9508_o;
  wire [63:0] n9509_o;
  wire n9510_o;
  wire n9511_o;
  wire [5:0] n9514_o;
  wire n9516_o;
  wire n9518_o;
  wire n9519_o;
  wire n9520_o;
  wire n9521_o;
  wire n9522_o;
  wire n9523_o;
  wire n9524_o;
  wire n9525_o;
  wire n9526_o;
  wire n9527_o;
  wire n9528_o;
  wire n9529_o;
  wire n9530_o;
  wire n9531_o;
  wire n9532_o;
  wire n9533_o;
  wire n9534_o;
  wire n9535_o;
  wire n9536_o;
  wire n9537_o;
  wire n9538_o;
  wire n9539_o;
  wire n9540_o;
  wire n9541_o;
  wire n9542_o;
  wire n9543_o;
  wire n9544_o;
  wire n9545_o;
  wire n9546_o;
  wire n9547_o;
  wire n9548_o;
  wire n9549_o;
  wire n9550_o;
  wire n9551_o;
  wire n9552_o;
  wire n9553_o;
  wire n9554_o;
  wire n9555_o;
  wire n9556_o;
  wire n9557_o;
  wire n9558_o;
  wire n9559_o;
  wire n9560_o;
  wire n9561_o;
  wire n9562_o;
  wire n9563_o;
  wire n9564_o;
  wire n9565_o;
  wire n9566_o;
  wire n9567_o;
  wire n9568_o;
  wire n9569_o;
  wire n9570_o;
  wire n9571_o;
  wire n9572_o;
  wire n9573_o;
  wire n9574_o;
  wire n9575_o;
  wire n9576_o;
  wire n9577_o;
  wire n9578_o;
  wire n9579_o;
  wire n9580_o;
  wire n9581_o;
  wire n9582_o;
  wire n9583_o;
  wire n9584_o;
  wire n9585_o;
  wire [3:0] n9586_o;
  wire [3:0] n9587_o;
  wire [3:0] n9588_o;
  wire [3:0] n9589_o;
  wire [3:0] n9590_o;
  wire [3:0] n9591_o;
  wire [3:0] n9592_o;
  wire [3:0] n9593_o;
  wire [3:0] n9594_o;
  wire [3:0] n9595_o;
  wire [3:0] n9596_o;
  wire [3:0] n9597_o;
  wire [3:0] n9598_o;
  wire [3:0] n9599_o;
  wire [3:0] n9600_o;
  wire [3:0] n9601_o;
  wire [15:0] n9602_o;
  wire [15:0] n9603_o;
  wire [15:0] n9604_o;
  wire [15:0] n9605_o;
  wire [63:0] n9606_o;
  wire [63:0] n9608_o;
  wire [127:0] n9609_o;
  wire [127:0] n9611_o;
  wire n9613_o;
  wire [127:0] n9614_o;
  wire [127:0] n9615_o;
  wire n9616_o;
  wire n9617_o;
  wire n9618_o;
  wire n9619_o;
  wire n9620_o;
  wire n9621_o;
  wire n9622_o;
  wire n9623_o;
  wire [5:0] n9624_o;
  wire n9626_o;
  wire n9628_o;
  wire [31:0] n9629_o;
  wire [63:0] n9631_o;
  wire [31:0] n9632_o;
  wire [63:0] n9634_o;
  wire [5:0] n9636_o;
  wire n9638_o;
  wire [31:0] n9639_o;
  wire [63:0] n9641_o;
  wire [31:0] n9642_o;
  wire [63:0] n9644_o;
  wire [63:0] n9645_o;
  wire [31:0] n9646_o;
  wire [63:0] n9648_o;
  wire [127:0] n9649_o;
  wire [127:0] n9650_o;
  wire [127:0] n9651_o;
  wire [127:0] n9652_o;
  wire [127:0] n9653_o;
  wire [127:0] n9654_o;
  wire n9655_o;
  wire [1:0] n9656_o;
  wire [63:0] n9657_o;
  wire n9659_o;
  wire [63:0] n9660_o;
  wire n9662_o;
  wire [31:0] n9663_o;
  wire [31:0] n9664_o;
  wire [63:0] n9665_o;
  wire n9667_o;
  wire [63:0] n9668_o;
  wire [2:0] n9669_o;
  reg [63:0] n9670_o;
  wire [2:0] n9671_o;
  wire n9673_o;
  wire n9674_o;
  wire n9675_o;
  wire n9676_o;
  wire n9677_o;
  wire n9678_o;
  wire n9679_o;
  wire [3:0] n9682_o;
  localparam [63:0] n9683_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire n9685_o;
  wire n9686_o;
  wire n9687_o;
  wire n9688_o;
  wire n9689_o;
  wire n9690_o;
  wire [3:0] n9692_o;
  wire [3:0] n9693_o;
  wire n9695_o;
  wire n9696_o;
  wire n9697_o;
  wire n9698_o;
  wire n9699_o;
  wire n9700_o;
  wire [3:0] n9702_o;
  wire [3:0] n9703_o;
  wire n9705_o;
  wire n9706_o;
  wire n9707_o;
  wire n9708_o;
  wire n9709_o;
  wire n9710_o;
  wire [3:0] n9712_o;
  wire [3:0] n9713_o;
  wire n9715_o;
  wire n9716_o;
  wire n9717_o;
  wire n9718_o;
  wire n9719_o;
  wire n9720_o;
  wire [3:0] n9722_o;
  wire [3:0] n9723_o;
  wire n9725_o;
  wire n9726_o;
  wire n9727_o;
  wire n9728_o;
  wire n9729_o;
  wire n9730_o;
  wire [3:0] n9732_o;
  wire [3:0] n9733_o;
  wire n9735_o;
  wire n9736_o;
  wire n9737_o;
  wire n9738_o;
  wire n9739_o;
  wire n9740_o;
  wire [3:0] n9742_o;
  wire [3:0] n9743_o;
  wire n9745_o;
  wire n9746_o;
  wire n9747_o;
  wire n9748_o;
  wire n9749_o;
  wire n9750_o;
  wire [3:0] n9752_o;
  wire [3:0] n9753_o;
  wire n9755_o;
  wire n9756_o;
  wire n9757_o;
  wire n9758_o;
  wire n9759_o;
  wire n9760_o;
  wire [3:0] n9762_o;
  wire [3:0] n9763_o;
  wire n9765_o;
  wire n9766_o;
  wire n9767_o;
  wire n9768_o;
  wire n9769_o;
  wire n9770_o;
  wire [3:0] n9772_o;
  wire [3:0] n9773_o;
  wire n9775_o;
  wire n9776_o;
  wire n9777_o;
  wire n9778_o;
  wire n9779_o;
  wire n9780_o;
  wire [3:0] n9782_o;
  wire [3:0] n9783_o;
  wire n9785_o;
  wire n9786_o;
  wire n9787_o;
  wire n9788_o;
  wire n9789_o;
  wire n9790_o;
  wire [3:0] n9792_o;
  wire [3:0] n9793_o;
  wire n9795_o;
  wire n9796_o;
  wire n9797_o;
  wire n9798_o;
  wire n9799_o;
  wire n9800_o;
  wire [3:0] n9802_o;
  wire [3:0] n9803_o;
  wire n9805_o;
  wire n9806_o;
  wire n9807_o;
  wire n9808_o;
  wire n9809_o;
  wire n9810_o;
  wire [3:0] n9812_o;
  wire [3:0] n9813_o;
  wire n9815_o;
  wire n9816_o;
  wire n9817_o;
  wire n9818_o;
  wire n9819_o;
  wire n9820_o;
  wire [3:0] n9822_o;
  wire [3:0] n9823_o;
  wire [3:0] n9824_o;
  wire n9825_o;
  wire n9826_o;
  wire [3:0] n9828_o;
  wire [63:0] n9829_o;
  wire n9831_o;
  wire [31:0] n9833_o;
  wire [4:0] n9838_o;
  wire [31:0] n9840_o;
  wire [31:0] n9842_o;
  wire [4:0] n9843_o;
  wire [63:0] n9846_o;
  wire n9848_o;
  wire n9849_o;
  wire [1:0] n9850_o;
  wire [31:0] n9851_o;
  wire [63:0] n9853_o;
  wire n9855_o;
  wire n9857_o;
  wire [1:0] n9858_o;
  reg [63:0] n9859_o;
  wire [63:0] n9861_o;
  wire n9864_o;
  wire [63:0] n9865_o;
  wire n9867_o;
  wire n9868_o;
  wire n9869_o;
  wire [63:0] n9871_o;
  wire [31:0] n9874_o;
  wire [7:0] n9879_o;
  wire n9884_o;
  wire n9888_o;
  wire n9892_o;
  wire [2:0] n9894_o;
  wire n9895_o;
  wire n9898_o;
  wire n9900_o;
  wire [2:0] n9901_o;
  wire n9902_o;
  wire n9903_o;
  wire n9904_o;
  wire n9905_o;
  wire n9906_o;
  wire n9907_o;
  wire n9908_o;
  wire n9911_o;
  wire n9913_o;
  wire [2:0] n9914_o;
  wire n9915_o;
  wire n9916_o;
  wire n9917_o;
  wire n9918_o;
  wire n9919_o;
  wire n9920_o;
  wire n9921_o;
  wire n9924_o;
  wire n9926_o;
  wire [2:0] n9927_o;
  wire n9928_o;
  wire n9929_o;
  wire n9930_o;
  wire n9931_o;
  wire n9932_o;
  wire n9933_o;
  wire n9934_o;
  wire n9937_o;
  wire n9939_o;
  wire [2:0] n9940_o;
  wire n9941_o;
  wire n9942_o;
  wire n9943_o;
  wire n9944_o;
  wire n9945_o;
  wire n9946_o;
  wire n9947_o;
  wire n9950_o;
  wire n9952_o;
  wire [2:0] n9953_o;
  wire n9954_o;
  wire n9955_o;
  wire n9956_o;
  wire n9957_o;
  wire n9958_o;
  wire n9959_o;
  wire n9960_o;
  wire n9963_o;
  wire n9965_o;
  wire [2:0] n9966_o;
  wire n9967_o;
  wire n9968_o;
  wire n9969_o;
  wire n9970_o;
  wire n9971_o;
  wire n9972_o;
  wire n9973_o;
  wire n9978_o;
  wire [2:0] n9979_o;
  wire n9981_o;
  wire n9982_o;
  wire n9984_o;
  wire n9985_o;
  wire [2:0] n9991_o;
  wire [31:0] n9992_o;
  wire n9994_o;
  wire [3:0] n9995_o;
  wire [3:0] n9997_o;
  localparam [63:0] n9998_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] n9999_o;
  wire [31:0] n10001_o;
  wire n10003_o;
  wire [3:0] n10004_o;
  wire [3:0] n10005_o;
  wire [3:0] n10006_o;
  wire [31:0] n10008_o;
  wire n10010_o;
  wire [3:0] n10011_o;
  wire [3:0] n10012_o;
  wire [3:0] n10013_o;
  wire [31:0] n10015_o;
  wire n10017_o;
  wire [3:0] n10018_o;
  wire [3:0] n10019_o;
  wire [3:0] n10020_o;
  wire [31:0] n10022_o;
  wire n10024_o;
  wire [3:0] n10025_o;
  wire [3:0] n10026_o;
  wire [3:0] n10027_o;
  wire [31:0] n10029_o;
  wire n10031_o;
  wire [3:0] n10032_o;
  wire [3:0] n10033_o;
  wire [3:0] n10034_o;
  wire [31:0] n10036_o;
  wire n10038_o;
  wire [3:0] n10039_o;
  wire [3:0] n10040_o;
  wire [3:0] n10041_o;
  wire [3:0] n10042_o;
  wire [31:0] n10043_o;
  wire n10045_o;
  wire [3:0] n10046_o;
  wire [3:0] n10047_o;
  wire [63:0] n10048_o;
  wire [63:0] n10049_o;
  wire n10056_o;
  wire [31:0] n10058_o;
  wire [2:0] n10063_o;
  wire [30:0] n10064_o;
  wire [31:0] n10065_o;
  wire [31:0] n10067_o;
  wire [4:0] n10068_o;
  wire [31:0] n10069_o;
  wire [31:0] n10071_o;
  wire [4:0] n10072_o;
  wire [31:0] n10075_o;
  wire [31:0] n10077_o;
  wire [4:0] n10078_o;
  wire n10083_o;
  wire n10085_o;
  wire [62:0] n10088_o;
  wire [63:0] n10091_o;
  wire n10093_o;
  wire [6:0] n10094_o;
  reg [63:0] n10097_o;
  wire [5:0] n10144_o;
  wire n10146_o;
  wire [31:0] n10148_o;
  wire n10153_o;
  wire n10154_o;
  wire n10155_o;
  wire n10156_o;
  wire [31:0] n10157_o;
  wire [31:0] n10158_o;
  wire [31:0] n10159_o;
  wire n10160_o;
  wire n10161_o;
  wire [31:0] n10162_o;
  wire [31:0] n10163_o;
  wire [31:0] n10164_o;
  wire n10165_o;
  wire n10166_o;
  wire n10167_o;
  wire n10168_o;
  wire n10169_o;
  wire [30:0] n10170_o;
  wire [30:0] n10171_o;
  wire n10172_o;
  wire n10175_o;
  wire [31:0] n10177_o;
  wire [31:0] n10178_o;
  wire n10179_o;
  wire n10182_o;
  wire n10184_o;
  wire n10185_o;
  wire n10186_o;
  wire n10187_o;
  wire n10188_o;
  wire n10189_o;
  wire n10190_o;
  wire n10191_o;
  wire n10192_o;
  wire n10193_o;
  wire n10194_o;
  wire n10195_o;
  wire n10196_o;
  wire n10197_o;
  wire [1:0] n10198_o;
  wire [2:0] n10200_o;
  wire [3:0] n10201_o;
  wire [4:0] n10202_o;
  wire n10203_o;
  wire [1:0] n10204_o;
  wire [2:0] n10206_o;
  wire [3:0] n10207_o;
  wire n10208_o;
  wire [4:0] n10209_o;
  wire [4:0] n10210_o;
  wire [4:0] n10212_o;
  wire [31:0] n10219_o;
  wire [2:0] n10224_o;
  wire [2:0] n10226_o;
  wire n10227_o;
  wire [2:0] n10228_o;
  wire n10229_o;
  wire [3:0] n10230_o;
  wire [1:0] n10231_o;
  wire n10232_o;
  wire [2:0] n10233_o;
  wire n10234_o;
  wire [3:0] n10235_o;
  wire [3:0] n10236_o;
  wire n10238_o;
  wire [31:0] n10241_o;
  wire n10246_o;
  wire [7:0] n10253_o;
  wire [7:0] n10255_o;
  wire n10256_o;
  wire [7:0] n10257_o;
  wire n10258_o;
  wire n10259_o;
  wire [7:0] n10260_o;
  wire n10261_o;
  wire n10262_o;
  wire [7:0] n10263_o;
  wire n10264_o;
  wire n10265_o;
  wire n10268_o;
  wire n10270_o;
  wire [1:0] n10273_o;
  wire [3:0] n10275_o;
  wire n10277_o;
  wire [7:0] n10285_o;
  wire [7:0] n10286_o;
  wire n10287_o;
  wire n10290_o;
  wire [7:0] n10292_o;
  wire [7:0] n10293_o;
  wire n10294_o;
  wire n10296_o;
  wire [7:0] n10297_o;
  wire [7:0] n10298_o;
  wire n10299_o;
  wire n10301_o;
  wire [7:0] n10302_o;
  wire [7:0] n10303_o;
  wire n10304_o;
  wire n10306_o;
  wire [7:0] n10307_o;
  wire [7:0] n10308_o;
  wire n10309_o;
  wire n10311_o;
  wire [7:0] n10312_o;
  wire [7:0] n10313_o;
  wire n10314_o;
  wire n10316_o;
  wire [7:0] n10317_o;
  wire [7:0] n10318_o;
  wire n10319_o;
  wire n10321_o;
  wire [7:0] n10322_o;
  wire [7:0] n10323_o;
  wire n10324_o;
  wire n10326_o;
  wire [1:0] n10328_o;
  wire [3:0] n10330_o;
  wire n10332_o;
  wire n10333_o;
  wire [2:0] n10342_o;
  wire [31:0] n10346_o;
  wire [4:0] n10351_o;
  wire [31:0] n10353_o;
  wire [4:0] n10358_o;
  wire [31:0] n10360_o;
  wire [4:0] n10365_o;
  wire [1:0] n10366_o;
  wire [30:0] n10367_o;
  wire [31:0] n10368_o;
  wire [31:0] n10370_o;
  wire [1:0] n10371_o;
  wire [30:0] n10372_o;
  wire [31:0] n10373_o;
  wire [31:0] n10375_o;
  wire [4:0] n10376_o;
  wire [30:0] n10377_o;
  wire [31:0] n10378_o;
  wire [31:0] n10380_o;
  wire [4:0] n10381_o;
  wire [1:0] n10386_o;
  wire [30:0] n10387_o;
  wire [31:0] n10388_o;
  wire [31:0] n10390_o;
  wire [4:0] n10391_o;
  wire [31:0] n10394_o;
  wire n10396_o;
  wire n10397_o;
  wire n10398_o;
  wire [31:0] n10400_o;
  wire n10402_o;
  wire n10403_o;
  wire n10404_o;
  wire [31:0] n10406_o;
  wire n10408_o;
  wire n10409_o;
  wire n10410_o;
  wire n10411_o;
  wire [31:0] n10412_o;
  wire n10414_o;
  wire n10415_o;
  wire [31:0] n10417_o;
  wire [2:0] n10422_o;
  wire [2:0] n10432_o;
  wire [3:0] n10435_o;
  wire [3:0] n10436_o;
  wire n10449_o;
  wire n10450_o;
  wire n10451_o;
  wire [1:0] n10452_o;
  wire n10453_o;
  wire [2:0] n10454_o;
  wire n10455_o;
  wire [3:0] n10456_o;
  wire n10458_o;
  wire [4:0] n10459_o;
  reg [3:0] n10461_o;
  wire [5:0] n10474_o;
  wire n10476_o;
  wire n10477_o;
  wire n10478_o;
  wire [31:0] n10480_o;
  wire [7:0] n10485_o;
  wire [31:0] n10488_o;
  wire [7:0] n10493_o;
  wire n10498_o;
  wire n10502_o;
  wire n10506_o;
  wire [2:0] n10508_o;
  wire n10509_o;
  wire n10512_o;
  wire n10514_o;
  wire [2:0] n10515_o;
  wire n10516_o;
  wire n10517_o;
  wire n10518_o;
  wire n10519_o;
  wire n10520_o;
  wire n10521_o;
  wire n10522_o;
  wire n10525_o;
  wire n10527_o;
  wire [2:0] n10528_o;
  wire n10529_o;
  wire n10530_o;
  wire n10531_o;
  wire n10532_o;
  wire n10533_o;
  wire n10534_o;
  wire n10535_o;
  wire n10538_o;
  wire n10540_o;
  wire [2:0] n10541_o;
  wire n10542_o;
  wire n10543_o;
  wire n10544_o;
  wire n10545_o;
  wire n10546_o;
  wire n10547_o;
  wire n10548_o;
  wire n10551_o;
  wire n10553_o;
  wire [2:0] n10554_o;
  wire n10555_o;
  wire n10556_o;
  wire n10557_o;
  wire n10558_o;
  wire n10559_o;
  wire n10560_o;
  wire n10561_o;
  wire n10564_o;
  wire n10566_o;
  wire [2:0] n10567_o;
  wire n10568_o;
  wire n10569_o;
  wire n10570_o;
  wire n10571_o;
  wire n10572_o;
  wire n10573_o;
  wire n10574_o;
  wire n10577_o;
  wire n10579_o;
  wire [2:0] n10580_o;
  wire n10581_o;
  wire n10582_o;
  wire n10583_o;
  wire n10584_o;
  wire n10585_o;
  wire n10586_o;
  wire n10587_o;
  wire n10592_o;
  wire [2:0] n10593_o;
  wire n10595_o;
  wire n10596_o;
  wire n10598_o;
  wire n10599_o;
  wire [2:0] n10605_o;
  wire n10613_o;
  wire n10616_o;
  wire n10619_o;
  wire n10622_o;
  wire n10625_o;
  wire n10628_o;
  wire n10631_o;
  wire n10634_o;
  wire [7:0] n10636_o;
  reg [7:0] n10637_o;
  wire [7:0] n10638_o;
  wire [31:0] n10640_o;
  wire n10648_o;
  wire n10651_o;
  wire n10654_o;
  wire n10657_o;
  wire n10660_o;
  wire n10663_o;
  wire n10666_o;
  wire n10669_o;
  wire [7:0] n10671_o;
  reg [7:0] n10672_o;
  wire [7:0] n10673_o;
  wire [11:0] n10674_o;
  wire [15:0] n10675_o;
  wire [19:0] n10676_o;
  wire [23:0] n10677_o;
  wire [27:0] n10678_o;
  wire [31:0] n10679_o;
  wire [7:0] n10680_o;
  wire [31:0] n10681_o;
  localparam [353:0] n10704_o = 354'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire n10706_o;
  wire n10707_o;
  wire n10708_o;
  wire [1:0] n10709_o;
  wire n10710_o;
  wire n10711_o;
  wire [2:0] n10712_o;
  wire n10713_o;
  wire n10714_o;
  wire [3:0] n10715_o;
  wire [31:0] n10737_o;
  wire n10740_o;
  wire n10741_o;
  wire n10742_o;
  wire n10743_o;
  wire n10744_o;
  wire n10745_o;
  wire [63:0] n10746_o;
  wire [63:0] n10748_o;
  wire [63:0] n10750_o;
  wire [63:0] n10752_o;
  wire [127:0] n10753_o;
  wire n10754_o;
  wire n10755_o;
  wire n10756_o;
  wire n10757_o;
  wire n10758_o;
  wire n10759_o;
  wire [391:0] n10764_o;
  wire [63:0] n10765_o;
  wire [63:0] n10767_o;
  wire [5:0] n10769_o;
  wire n10771_o;
  wire n10772_o;
  wire [5:0] n10775_o;
  wire n10777_o;
  wire [5:0] n10778_o;
  wire n10780_o;
  wire n10781_o;
  wire n10782_o;
  wire [5:0] n10785_o;
  wire n10787_o;
  wire [5:0] n10788_o;
  wire n10790_o;
  wire n10791_o;
  wire n10792_o;
  wire [5:0] n10795_o;
  wire n10797_o;
  wire n10798_o;
  wire [5:0] n10801_o;
  wire n10803_o;
  wire n10804_o;
  wire n10806_o;
  wire [353:0] n10809_o;
  wire [11:0] n10810_o;
  wire [11:0] n10811_o;
  wire [11:0] n10812_o;
  wire n10815_o;
  wire n10816_o;
  wire [63:0] n10817_o;
  wire [63:0] n10819_o;
  wire [353:0] n10820_o;
  wire [63:0] n10821_o;
  wire [63:0] n10822_o;
  wire [66:0] n10823_o;
  wire n10824_o;
  wire n10825_o;
  wire [113:0] n10826_o;
  wire [2:0] n10828_o;
  wire n10829_o;
  wire n10830_o;
  wire n10831_o;
  wire n10832_o;
  wire [5:0] n10833_o;
  wire [391:0] n10834_o;
  wire [5:0] n10835_o;
  wire [5:0] n10836_o;
  wire n10837_o;
  wire n10839_o;
  wire n10840_o;
  wire n10841_o;
  wire n10842_o;
  wire n10843_o;
  wire n10844_o;
  wire n10845_o;
  wire n10846_o;
  wire n10848_o;
  wire n10852_o;
  wire [5:0] n10855_o;
  wire n10857_o;
  wire [5:0] n10858_o;
  wire n10860_o;
  wire n10861_o;
  wire [5:0] n10862_o;
  wire n10864_o;
  wire n10865_o;
  wire [5:0] n10866_o;
  wire n10868_o;
  wire n10869_o;
  wire [5:0] n10870_o;
  wire n10872_o;
  wire n10873_o;
  wire [5:0] n10874_o;
  wire n10876_o;
  wire n10877_o;
  wire [5:0] n10879_o;
  wire n10881_o;
  wire [5:0] n10882_o;
  wire n10884_o;
  wire n10885_o;
  wire [5:0] n10886_o;
  wire n10888_o;
  wire n10889_o;
  wire n10891_o;
  wire n10892_o;
  wire n10893_o;
  wire n10894_o;
  wire n10895_o;
  wire n10896_o;
  wire n10897_o;
  wire n10898_o;
  wire n10899_o;
  wire n10900_o;
  wire n10901_o;
  wire n10902_o;
  wire n10903_o;
  wire n10905_o;
  wire [11:0] n10909_o;
  wire n10910_o;
  wire [11:0] n10911_o;
  wire n10912_o;
  wire [11:0] n10913_o;
  wire n10914_o;
  wire n10915_o;
  wire [5:0] n10917_o;
  wire [31:0] n10918_o;
  wire [5:0] n10924_o;
  wire n10929_o;
  wire n10932_o;
  wire n10934_o;
  wire n10935_o;
  wire n10936_o;
  wire n10938_o;
  wire n10939_o;
  wire n10940_o;
  wire n10943_o;
  wire n10944_o;
  wire n10946_o;
  wire n10947_o;
  wire n10949_o;
  wire n10950_o;
  wire [11:0] n10952_o;
  wire n10954_o;
  wire [11:0] n10955_o;
  wire n10956_o;
  wire n10957_o;
  wire n10958_o;
  wire n10959_o;
  wire n10961_o;
  wire [11:0] n10962_o;
  wire n10963_o;
  wire n10964_o;
  wire n10965_o;
  wire n10966_o;
  wire n10967_o;
  wire n10969_o;
  wire [1:0] n10970_o;
  wire [11:0] n10971_o;
  wire n10972_o;
  wire n10973_o;
  wire n10974_o;
  wire n10975_o;
  wire [1:0] n10976_o;
  wire [1:0] n10977_o;
  wire [1:0] n10978_o;
  wire [1:0] n10979_o;
  wire n10980_o;
  wire n10981_o;
  wire n10982_o;
  wire n10983_o;
  wire n10984_o;
  wire n10986_o;
  wire [11:0] n10987_o;
  wire n10988_o;
  wire n10989_o;
  wire n10990_o;
  wire n10991_o;
  wire n10992_o;
  wire n10993_o;
  wire n10994_o;
  wire n10995_o;
  wire n10996_o;
  wire n10997_o;
  wire n10998_o;
  wire n10999_o;
  wire [1:0] n11000_o;
  wire [1:0] n11001_o;
  wire [1:0] n11002_o;
  wire [1:0] n11003_o;
  wire n11004_o;
  wire n11005_o;
  wire n11006_o;
  wire n11007_o;
  wire n11008_o;
  wire n11010_o;
  wire [11:0] n11011_o;
  wire n11012_o;
  wire n11013_o;
  wire n11014_o;
  wire n11015_o;
  wire n11016_o;
  wire n11017_o;
  wire n11018_o;
  wire n11019_o;
  wire n11020_o;
  wire n11021_o;
  wire n11022_o;
  wire n11023_o;
  wire [1:0] n11024_o;
  wire [1:0] n11025_o;
  wire [1:0] n11026_o;
  wire [1:0] n11027_o;
  wire n11028_o;
  wire n11029_o;
  wire n11030_o;
  wire n11031_o;
  wire n11032_o;
  wire n11039_o;
  wire n11040_o;
  wire n11041_o;
  wire n11045_o;
  wire n11046_o;
  wire n11047_o;
  wire [5:0] n11051_o;
  wire [5:0] n11052_o;
  wire [5:0] n11053_o;
  wire n11054_o;
  wire n11055_o;
  wire n11056_o;
  wire n11057_o;
  wire n11058_o;
  wire n11059_o;
  wire n11060_o;
  wire n11061_o;
  wire n11062_o;
  wire n11065_o;
  wire n11066_o;
  wire n11067_o;
  wire [1:0] n11068_o;
  wire n11069_o;
  wire n11071_o;
  wire n11072_o;
  wire n11073_o;
  wire n11074_o;
  wire n11075_o;
  wire n11076_o;
  wire n11077_o;
  wire n11078_o;
  wire n11079_o;
  wire n11080_o;
  wire n11081_o;
  wire n11083_o;
  wire n11084_o;
  wire n11086_o;
  wire n11087_o;
  wire n11088_o;
  wire n11090_o;
  wire [1:0] n11091_o;
  wire n11093_o;
  wire n11094_o;
  wire [5:0] n11096_o;
  wire n11098_o;
  wire n11099_o;
  wire [11:0] n11101_o;
  wire [63:0] n11102_o;
  wire n11104_o;
  wire n11107_o;
  wire n11109_o;
  wire [9:0] n11110_o;
  wire n11112_o;
  wire n11114_o;
  wire n11117_o;
  wire n11119_o;
  wire n11121_o;
  wire n11123_o;
  wire n11124_o;
  wire n11126_o;
  wire n11127_o;
  wire n11129_o;
  wire n11130_o;
  wire n11132_o;
  wire n11133_o;
  wire n11135_o;
  wire n11136_o;
  wire n11137_o;
  wire [1:0] n11138_o;
  wire n11140_o;
  wire [798:0] n11142_o;
  wire [119:0] n11146_o;
  wire [231:0] n11147_o;
  wire [353:0] n11148_o;
  wire [1:0] n11149_o;
  wire [121:0] n11150_o;
  wire [1:0] n11151_o;
  wire [121:0] n11152_o;
  wire [121:0] n11153_o;
  wire [1:0] n11154_o;
  wire [1:0] n11155_o;
  wire [229:0] n11156_o;
  wire n11157_o;
  wire [229:0] n11158_o;
  wire [229:0] n11159_o;
  wire [353:0] n11160_o;
  wire [353:0] n11161_o;
  wire [353:0] n11162_o;
  wire n11163_o;
  wire [798:0] n11165_o;
  wire n11170_o;
  wire n11171_o;
  wire [121:0] n11172_o;
  wire [228:0] n11173_o;
  wire [353:0] n11174_o;
  wire [353:0] n11175_o;
  wire n11177_o;
  wire n11179_o;
  wire [31:0] n11183_o;
  wire [4:0] n11188_o;
  wire [4:0] n11189_o;
  wire n11190_o;
  wire n11192_o;
  wire n11194_o;
  wire n11196_o;
  wire n11198_o;
  wire n11200_o;
  wire n11202_o;
  wire n11204_o;
  wire n11205_o;
  wire n11207_o;
  wire n11208_o;
  wire n11210_o;
  wire n11211_o;
  wire n11213_o;
  wire n11214_o;
  wire n11216_o;
  wire n11217_o;
  wire n11219_o;
  wire n11220_o;
  wire n11222_o;
  wire n11223_o;
  wire n11224_o;
  wire n11225_o;
  wire n11227_o;
  wire n11230_o;
  wire [31:0] n11232_o;
  wire [4:0] n11237_o;
  wire [31:0] n11239_o;
  wire [4:0] n11244_o;
  wire n11245_o;
  wire n11246_o;
  wire [30:0] n11257_o;
  wire [31:0] n11258_o;
  wire [31:0] n11261_o;
  wire [4:0] n11262_o;
  wire n11265_o;
  wire n11266_o;
  wire n11268_o;
  wire n11272_o;
  wire n11274_o;
  wire n11277_o;
  wire n11278_o;
  wire n11279_o;
  wire n11280_o;
  wire n11282_o;
  wire n11283_o;
  wire n11285_o;
  wire n11286_o;
  wire n11287_o;
  wire n11288_o;
  wire n11289_o;
  wire n11290_o;
  wire n11291_o;
  wire n11292_o;
  wire [5:0] n11293_o;
  wire n11295_o;
  wire n11298_o;
  wire n11299_o;
  wire n11301_o;
  wire n11304_o;
  wire n11306_o;
  wire n11307_o;
  wire n11309_o;
  wire n11311_o;
  wire n11312_o;
  wire n11313_o;
  wire n11314_o;
  wire n11315_o;
  wire n11316_o;
  wire n11317_o;
  wire [1:0] n11318_o;
  wire n11319_o;
  wire n11320_o;
  wire [2:0] n11321_o;
  wire n11322_o;
  wire n11323_o;
  wire [3:0] n11324_o;
  wire [32:0] n11325_o;
  wire [4:0] n11326_o;
  wire n11328_o;
  wire [1:0] n11332_o;
  wire [1:0] n11333_o;
  wire [1:0] n11334_o;
  wire n11335_o;
  wire n11336_o;
  wire [3:0] n11338_o;
  wire [8:0] n11339_o;
  wire n11340_o;
  wire n11341_o;
  wire n11342_o;
  wire n11343_o;
  wire n11344_o;
  wire n11346_o;
  wire n11351_o;
  wire n11353_o;
  wire n11354_o;
  wire n11356_o;
  wire n11358_o;
  wire n11360_o;
  wire n11362_o;
  wire n11364_o;
  wire [6:0] n11366_o;
  wire n11371_o;
  wire [31:0] n11373_o;
  wire [4:0] n11378_o;
  wire [4:0] n11379_o;
  wire [9:0] n11380_o;
  wire [31:0] n11382_o;
  wire n11384_o;
  wire n11386_o;
  wire n11387_o;
  wire n11388_o;
  wire n11390_o;
  wire n11391_o;
  wire [45:0] n11392_o;
  wire [45:0] n11393_o;
  wire [45:0] n11394_o;
  wire [17:0] n11395_o;
  wire [31:0] n11397_o;
  wire [4:0] n11402_o;
  wire [4:0] n11403_o;
  wire [9:0] n11404_o;
  wire [63:0] n11406_o;
  wire n11408_o;
  wire [31:0] n11410_o;
  wire n11412_o;
  wire [63:0] n11413_o;
  wire n11415_o;
  wire [63:0] n11416_o;
  wire n11418_o;
  wire n11422_o;
  wire [31:0] n11423_o;
  wire [63:0] n11424_o;
  wire n11426_o;
  wire [31:0] n11427_o;
  wire [31:0] n11429_o;
  wire n11431_o;
  wire [63:0] n11433_o;
  wire n11435_o;
  wire n11437_o;
  wire n11438_o;
  wire n11440_o;
  wire n11441_o;
  wire n11443_o;
  wire n11444_o;
  wire n11446_o;
  wire n11447_o;
  wire n11449_o;
  wire n11450_o;
  wire n11452_o;
  wire n11453_o;
  wire n11455_o;
  wire n11456_o;
  wire n11458_o;
  wire n11459_o;
  wire n11461_o;
  wire n11462_o;
  wire n11464_o;
  wire n11465_o;
  wire n11467_o;
  wire n11468_o;
  wire n11470_o;
  wire n11471_o;
  wire n11473_o;
  wire n11474_o;
  wire n11476_o;
  wire n11477_o;
  wire n11479_o;
  wire n11480_o;
  wire n11482_o;
  wire n11483_o;
  wire n11485_o;
  wire n11486_o;
  wire n11488_o;
  wire n11489_o;
  wire n11491_o;
  wire n11492_o;
  wire n11494_o;
  wire n11495_o;
  wire n11497_o;
  wire n11498_o;
  wire n11500_o;
  wire n11501_o;
  wire n11503_o;
  wire n11504_o;
  wire n11506_o;
  wire n11507_o;
  wire n11509_o;
  wire n11510_o;
  wire [6:0] n11512_o;
  wire n11517_o;
  wire n11518_o;
  wire n11519_o;
  wire n11520_o;
  wire n11523_o;
  wire [7:0] n11524_o;
  reg n11525_o;
  reg [31:0] n11526_o;
  reg n11528_o;
  wire [31:0] n11529_o;
  wire [31:0] n11530_o;
  wire [31:0] n11531_o;
  wire [31:0] n11532_o;
  wire [31:0] n11533_o;
  wire [31:0] n11534_o;
  wire [31:0] n11535_o;
  reg [31:0] n11536_o;
  wire [31:0] n11537_o;
  wire [31:0] n11538_o;
  wire [31:0] n11539_o;
  wire [31:0] n11540_o;
  wire [31:0] n11541_o;
  wire [31:0] n11542_o;
  wire [31:0] n11543_o;
  reg [31:0] n11544_o;
  wire n11546_o;
  wire [31:0] n11547_o;
  wire n11549_o;
  wire [63:0] n11550_o;
  wire [63:0] n11551_o;
  wire [63:0] n11552_o;
  wire n11554_o;
  wire n11556_o;
  wire n11558_o;
  wire n11559_o;
  wire n11560_o;
  wire n11561_o;
  wire n11562_o;
  wire n11563_o;
  wire [2:0] n11564_o;
  wire [27:0] n11565_o;
  wire [27:0] n11566_o;
  wire [27:0] n11567_o;
  wire [2:0] n11568_o;
  wire [2:0] n11569_o;
  wire n11572_o;
  wire [1:0] n11576_o;
  wire [1:0] n11577_o;
  wire [1:0] n11578_o;
  wire n11579_o;
  wire n11580_o;
  wire [5:0] n11581_o;
  wire [2:0] n11582_o;
  wire [15:0] n11583_o;
  wire [1:0] n11584_o;
  wire n11585_o;
  wire n11586_o;
  wire n11587_o;
  wire n11588_o;
  wire n11589_o;
  wire [10:0] n11590_o;
  wire [46:0] n11591_o;
  wire n11592_o;
  wire n11593_o;
  wire [9:0] n11594_o;
  wire [9:0] n11595_o;
  wire [9:0] n11596_o;
  wire [1:0] n11597_o;
  wire [1:0] n11598_o;
  wire [1:0] n11599_o;
  wire n11600_o;
  wire n11601_o;
  wire [43:0] n11602_o;
  wire [43:0] n11603_o;
  wire [43:0] n11604_o;
  wire [2:0] n11605_o;
  wire [2:0] n11606_o;
  wire n11607_o;
  wire n11608_o;
  wire n11610_o;
  wire [6:0] n11612_o;
  wire n11617_o;
  wire [31:0] n11619_o;
  wire [4:0] n11624_o;
  wire [4:0] n11625_o;
  wire [9:0] n11626_o;
  wire [31:0] n11628_o;
  wire n11630_o;
  wire n11631_o;
  wire n11632_o;
  wire n11633_o;
  wire n11634_o;
  wire n11635_o;
  wire [4:0] n11636_o;
  wire [4:0] n11637_o;
  wire [31:0] n11639_o;
  wire [4:0] n11644_o;
  wire [4:0] n11645_o;
  wire [9:0] n11646_o;
  wire n11649_o;
  wire [31:0] n11650_o;
  wire n11652_o;
  wire n11655_o;
  wire n11657_o;
  wire n11658_o;
  wire n11660_o;
  wire n11661_o;
  wire n11663_o;
  wire n11664_o;
  wire n11666_o;
  wire n11667_o;
  wire n11669_o;
  wire n11670_o;
  wire n11672_o;
  wire n11673_o;
  wire n11675_o;
  wire n11676_o;
  wire n11678_o;
  wire n11679_o;
  wire n11681_o;
  wire n11682_o;
  wire n11684_o;
  wire n11685_o;
  wire n11687_o;
  wire n11688_o;
  wire n11690_o;
  wire n11691_o;
  wire n11693_o;
  wire n11694_o;
  wire n11696_o;
  wire n11697_o;
  wire n11699_o;
  wire n11700_o;
  wire n11702_o;
  wire n11703_o;
  wire n11705_o;
  wire n11706_o;
  wire n11708_o;
  wire n11709_o;
  wire n11711_o;
  wire n11712_o;
  wire n11714_o;
  wire n11715_o;
  wire n11717_o;
  wire n11718_o;
  wire n11719_o;
  wire n11722_o;
  wire [2:0] n11723_o;
  reg [63:0] n11724_o;
  reg n11725_o;
  reg [31:0] n11726_o;
  reg n11728_o;
  wire [63:0] n11729_o;
  wire n11730_o;
  wire n11731_o;
  wire [31:0] n11732_o;
  wire n11734_o;
  wire n11736_o;
  wire n11737_o;
  wire [798:0] n11739_o;
  wire [119:0] n11743_o;
  wire [231:0] n11744_o;
  wire [353:0] n11745_o;
  wire [353:0] n11746_o;
  wire [353:0] n11747_o;
  wire n11749_o;
  wire n11751_o;
  wire n11752_o;
  wire n11754_o;
  wire n11755_o;
  wire n11757_o;
  wire n11758_o;
  wire n11760_o;
  wire n11761_o;
  wire n11763_o;
  wire n11764_o;
  wire n11766_o;
  wire n11770_o;
  wire n11772_o;
  wire n11778_o;
  wire n11780_o;
  wire n11781_o;
  wire n11783_o;
  wire n11784_o;
  wire n11790_o;
  wire n11792_o;
  wire n11793_o;
  wire n11795_o;
  wire n11796_o;
  wire [30:0] n11798_o;
  reg n11801_o;
  reg [63:0] n11802_o;
  wire n11803_o;
  wire n11804_o;
  reg n11805_o;
  wire n11806_o;
  wire n11807_o;
  reg n11808_o;
  wire [1:0] n11809_o;
  wire [1:0] n11810_o;
  wire [1:0] n11811_o;
  reg [1:0] n11812_o;
  wire [1:0] n11813_o;
  wire [1:0] n11814_o;
  reg [1:0] n11815_o;
  wire [5:0] n11816_o;
  wire [5:0] n11817_o;
  wire [5:0] n11818_o;
  reg [5:0] n11819_o;
  wire n11820_o;
  wire n11821_o;
  reg n11822_o;
  wire [1:0] n11823_o;
  wire [1:0] n11824_o;
  reg [1:0] n11825_o;
  wire n11826_o;
  reg n11827_o;
  wire [5:0] n11828_o;
  wire [5:0] n11829_o;
  reg [5:0] n11830_o;
  wire [4:0] n11831_o;
  wire [4:0] n11832_o;
  reg [4:0] n11833_o;
  wire [3:0] n11834_o;
  wire [3:0] n11835_o;
  reg [3:0] n11836_o;
  wire [28:0] n11837_o;
  wire [28:0] n11838_o;
  wire [28:0] n11839_o;
  reg [28:0] n11840_o;
  wire n11841_o;
  wire n11842_o;
  reg n11843_o;
  wire [2:0] n11844_o;
  wire [2:0] n11845_o;
  reg [2:0] n11846_o;
  reg [63:0] n11848_o;
  reg n11849_o;
  reg n11850_o;
  reg n11851_o;
  reg n11852_o;
  wire n11853_o;
  wire n11854_o;
  reg n11855_o;
  wire [118:0] n11856_o;
  wire [118:0] n11857_o;
  wire [118:0] n11858_o;
  reg [118:0] n11859_o;
  wire [4:0] n11860_o;
  wire [4:0] n11861_o;
  reg [4:0] n11862_o;
  wire n11863_o;
  wire n11864_o;
  reg n11865_o;
  wire [11:0] n11866_o;
  wire [11:0] n11867_o;
  reg [11:0] n11868_o;
  wire n11869_o;
  wire n11870_o;
  reg n11871_o;
  wire [3:0] n11872_o;
  wire [3:0] n11873_o;
  reg [3:0] n11874_o;
  wire [63:0] n11875_o;
  wire [63:0] n11876_o;
  reg [63:0] n11877_o;
  wire [63:0] n11878_o;
  wire [63:0] n11879_o;
  wire [63:0] n11880_o;
  reg [63:0] n11881_o;
  wire [3:0] n11882_o;
  wire [3:0] n11883_o;
  wire [2:0] n11884_o;
  wire [3:0] n11885_o;
  reg [3:0] n11886_o;
  wire n11887_o;
  wire n11888_o;
  reg n11889_o;
  wire [77:0] n11890_o;
  wire [77:0] n11891_o;
  wire [77:0] n11892_o;
  reg [77:0] n11893_o;
  reg n11894_o;
  reg n11895_o;
  wire n11896_o;
  reg n11897_o;
  reg n11898_o;
  reg n11899_o;
  reg n11900_o;
  reg n11901_o;
  reg n11902_o;
  reg [31:0] n11903_o;
  reg n11906_o;
  reg n11909_o;
  reg n11913_o;
  reg n11916_o;
  reg n11920_o;
  reg n11923_o;
  reg n11927_o;
  wire [63:0] n11928_o;
  wire [63:0] n11929_o;
  wire [63:0] n11930_o;
  wire [63:0] n11932_o;
  wire n11933_o;
  wire n11934_o;
  wire n11935_o;
  wire n11936_o;
  wire n11938_o;
  wire n11939_o;
  wire n11941_o;
  wire [66:0] n11942_o;
  wire n11943_o;
  wire [2:0] n11944_o;
  wire [66:0] n11945_o;
  wire [66:0] n11946_o;
  wire n11947_o;
  wire n11948_o;
  wire n11949_o;
  wire n11950_o;
  wire n11952_o;
  wire [1:0] n11953_o;
  wire n11955_o;
  wire [1:0] n11957_o;
  wire n11959_o;
  wire [1:0] n11960_o;
  wire n11962_o;
  wire n11964_o;
  wire n11967_o;
  wire n11970_o;
  wire n11972_o;
  wire n11974_o;
  wire n11976_o;
  wire n11978_o;
  wire [5:0] n11979_o;
  wire n11981_o;
  wire n11983_o;
  wire n11985_o;
  wire n11987_o;
  wire n11988_o;
  wire n11990_o;
  wire n11992_o;
  wire [191:0] n11994_o;
  wire [191:0] n11995_o;
  wire [63:0] n11998_o;
  wire n12000_o;
  wire n12001_o;
  wire [1:0] n12002_o;
  wire [1:0] n12003_o;
  wire [1:0] n12004_o;
  wire [353:0] n12005_o;
  wire [1:0] n12006_o;
  wire [1:0] n12007_o;
  wire [1:0] n12008_o;
  wire [33:0] n12009_o;
  wire [353:0] n12010_o;
  wire [1:0] n12012_o;
  wire n12014_o;
  wire n12015_o;
  wire [1:0] n12016_o;
  wire [1:0] n12018_o;
  wire [33:0] n12020_o;
  wire [33:0] n12021_o;
  wire n12022_o;
  wire n12026_o;
  localparam [389:0] n12027_o = 390'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire n12029_o;
  wire n12030_o;
  wire n12047_o;
  wire n12049_o;
  wire n12052_o;
  wire n12054_o;
  wire n12055_o;
  wire n12056_o;
  wire n12057_o;
  wire n12058_o;
  wire n12059_o;
  wire n12060_o;
  wire n12061_o;
  wire n12062_o;
  wire n12063_o;
  wire n12064_o;
  wire n12065_o;
  wire n12067_o;
  wire n12068_o;
  wire n12069_o;
  wire n12070_o;
  wire n12073_o;
  wire n12075_o;
  wire n12076_o;
  wire n12077_o;
  wire n12078_o;
  wire [2:0] n12079_o;
  wire [2:0] n12080_o;
  wire [2:0] n12081_o;
  wire [2:0] n12082_o;
  wire [2:0] n12083_o;
  wire n12085_o;
  wire n12086_o;
  wire n12087_o;
  wire n12088_o;
  wire [2:0] n12089_o;
  wire [2:0] n12090_o;
  wire [2:0] n12091_o;
  wire [2:0] n12092_o;
  wire n12093_o;
  wire n12094_o;
  wire n12095_o;
  wire n12096_o;
  wire n12097_o;
  wire n12099_o;
  wire n12100_o;
  wire n12101_o;
  wire n12102_o;
  wire n12103_o;
  wire n12104_o;
  wire [2:0] n12105_o;
  wire [2:0] n12106_o;
  wire [2:0] n12107_o;
  wire [2:0] n12108_o;
  wire n12109_o;
  wire n12110_o;
  wire n12111_o;
  wire n12112_o;
  wire n12113_o;
  wire n12114_o;
  wire n12115_o;
  wire n12116_o;
  wire n12117_o;
  wire n12118_o;
  wire n12120_o;
  wire n12121_o;
  wire n12122_o;
  wire n12123_o;
  wire n12125_o;
  wire n12126_o;
  wire n12127_o;
  wire n12128_o;
  wire [2:0] n12130_o;
  wire n12131_o;
  wire n12132_o;
  wire n12133_o;
  wire n12134_o;
  wire [2:0] n12135_o;
  wire [2:0] n12136_o;
  wire [2:0] n12137_o;
  wire [2:0] n12138_o;
  wire n12141_o;
  wire [2:0] n12142_o;
  wire n12143_o;
  wire [2:0] n12144_o;
  wire n12145_o;
  wire n12146_o;
  wire n12147_o;
  wire n12148_o;
  wire n12149_o;
  wire n12150_o;
  wire n12151_o;
  wire n12152_o;
  wire n12153_o;
  wire n12154_o;
  wire [2:0] n12155_o;
  wire [2:0] n12156_o;
  wire n12159_o;
  wire n12160_o;
  wire [2:0] n12161_o;
  wire [2:0] n12162_o;
  wire [2:0] n12163_o;
  wire [2:0] n12164_o;
  wire n12165_o;
  wire n12166_o;
  wire n12167_o;
  wire n12168_o;
  wire n12169_o;
  wire n12170_o;
  wire n12171_o;
  wire n12172_o;
  wire n12173_o;
  wire n12174_o;
  wire [2:0] n12175_o;
  wire [2:0] n12176_o;
  wire [120:0] n12183_o;
  wire [120:0] n12184_o;
  wire [120:0] n12185_o;
  wire n12186_o;
  wire n12187_o;
  wire n12188_o;
  wire n12189_o;
  wire n12190_o;
  wire n12191_o;
  wire n12192_o;
  wire n12193_o;
  wire n12194_o;
  wire n12197_o;
  wire [11:0] n12201_o;
  wire [11:0] n12202_o;
  wire [11:0] n12203_o;
  wire [11:0] n12204_o;
  wire n12205_o;
  wire n12206_o;
  wire n12207_o;
  wire n12208_o;
  wire [75:0] n12215_o;
  wire [75:0] n12216_o;
  wire [75:0] n12217_o;
  wire [138:0] n12218_o;
  wire [138:0] n12219_o;
  wire [138:0] n12220_o;
  wire n12222_o;
  wire n12223_o;
  wire n12224_o;
  wire n12225_o;
  wire n12226_o;
  wire n12227_o;
  wire [798:0] n12228_o;
  wire [353:0] n12229_o;
  wire n12230_o;
  wire n12232_o;
  wire n12234_o;
  wire [1:0] n12250_o;
  wire [1:0] n12251_o;
  wire [3:0] n12252_o;
  wire [2:0] n12253_o;
  wire [1:0] n12254_o;
  wire [1:0] n12255_o;
  wire [1:0] n12256_o;
  wire [1:0] n12257_o;
  wire [1:0] n12258_o;
  wire [1:0] n12259_o;
  wire [1:0] n12260_o;
  wire [1:0] n12261_o;
  wire [3:0] n12262_o;
  wire [3:0] n12263_o;
  wire [3:0] n12264_o;
  wire [3:0] n12265_o;
  wire [2:0] n12266_o;
  wire [2:0] n12267_o;
  wire [2:0] n12268_o;
  wire [2:0] n12269_o;
  wire n12270_o;
  wire n12271_o;
  wire n12272_o;
  wire n12273_o;
  wire [63:0] n12277_o;
  wire [63:0] n12278_o;
  wire [63:0] n12279_o;
  wire [1:0] n12283_o;
  wire [1:0] n12284_o;
  wire [1:0] n12285_o;
  wire [1:0] n12289_o;
  wire [1:0] n12290_o;
  wire [1:0] n12291_o;
  wire n12295_o;
  wire n12296_o;
  wire n12297_o;
  wire [63:0] n12298_o;
  wire [63:0] n12299_o;
  wire [63:0] n12300_o;
  wire [46:0] n12301_o;
  wire [46:0] n12302_o;
  wire [46:0] n12303_o;
  wire [2:0] n12304_o;
  wire [2:0] n12305_o;
  wire [2:0] n12306_o;
  wire n12307_o;
  wire [353:0] n12308_o;
  wire [63:0] n12309_o;
  wire [63:0] n12310_o;
  wire [43:0] n12311_o;
  wire [43:0] n12312_o;
  wire [43:0] n12313_o;
  wire [6:0] n12317_o;
  wire [5:0] n12318_o;
  wire [5:0] n12319_o;
  wire [5:0] n12320_o;
  wire n12321_o;
  wire [798:0] n12322_o;
  wire [353:0] n12323_o;
  wire n12324_o;
  wire n12325_o;
  wire n12326_o;
  wire n12327_o;
  wire [4:0] n12328_o;
  wire [4:0] n12329_o;
  wire [4:0] n12330_o;
  wire n12331_o;
  wire [798:0] n12332_o;
  wire [353:0] n12333_o;
  wire n12334_o;
  wire n12335_o;
  wire n12336_o;
  wire n12337_o;
  wire n12338_o;
  wire n12339_o;
  wire n12340_o;
  wire [2:0] n12341_o;
  wire [2:0] n12342_o;
  wire [2:0] n12343_o;
  wire [2:0] n12344_o;
  wire [2:0] n12345_o;
  wire [2:0] n12346_o;
  wire n12350_o;
  wire n12351_o;
  wire n12352_o;
  wire n12353_o;
  wire [798:0] n12354_o;
  wire [353:0] n12355_o;
  wire n12356_o;
  wire n12357_o;
  wire n12358_o;
  wire n12359_o;
  wire n12360_o;
  wire [798:0] n12361_o;
  wire [353:0] n12362_o;
  wire n12363_o;
  wire n12364_o;
  wire n12365_o;
  wire n12366_o;
  wire [1:0] n12367_o;
  wire [1:0] n12368_o;
  wire [1:0] n12369_o;
  wire [2:0] n12370_o;
  wire n12371_o;
  wire n12372_o;
  wire n12373_o;
  wire [798:0] n12374_o;
  wire [353:0] n12375_o;
  wire n12376_o;
  wire n12377_o;
  wire [2:0] n12378_o;
  wire [1:0] n12379_o;
  wire [798:0] n12380_o;
  wire [353:0] n12381_o;
  wire [63:0] n12382_o;
  wire [2:0] n12383_o;
  wire n12384_o;
  wire n12385_o;
  wire n12386_o;
  wire [798:0] n12387_o;
  wire [353:0] n12388_o;
  wire n12389_o;
  wire n12390_o;
  wire [2:0] n12391_o;
  wire [1:0] n12392_o;
  wire [798:0] n12393_o;
  wire n12394_o;
  wire [798:0] n12395_o;
  wire [3:0] n12396_o;
  wire [3:0] n12397_o;
  wire [3:0] n12398_o;
  wire [798:0] n12399_o;
  wire n12400_o;
  wire [798:0] n12401_o;
  wire [3:0] n12402_o;
  wire [3:0] n12403_o;
  wire [3:0] n12404_o;
  wire [798:0] n12405_o;
  wire n12406_o;
  wire [798:0] n12407_o;
  wire [3:0] n12408_o;
  wire [3:0] n12409_o;
  wire [3:0] n12410_o;
  wire [798:0] n12411_o;
  wire n12412_o;
  wire [798:0] n12413_o;
  wire [3:0] n12414_o;
  wire [3:0] n12415_o;
  wire [3:0] n12416_o;
  wire [798:0] n12417_o;
  wire n12418_o;
  wire [798:0] n12419_o;
  wire [3:0] n12420_o;
  wire [3:0] n12421_o;
  wire [3:0] n12422_o;
  wire [798:0] n12423_o;
  wire n12424_o;
  wire [798:0] n12425_o;
  wire [3:0] n12426_o;
  wire [3:0] n12427_o;
  wire [3:0] n12428_o;
  wire [798:0] n12429_o;
  wire n12430_o;
  wire [798:0] n12431_o;
  wire [3:0] n12432_o;
  wire [3:0] n12433_o;
  wire [3:0] n12434_o;
  wire [798:0] n12435_o;
  wire n12436_o;
  wire [798:0] n12437_o;
  wire [3:0] n12438_o;
  wire [3:0] n12439_o;
  wire [3:0] n12440_o;
  wire [5:0] n12441_o;
  wire [63:0] n12443_o;
  wire [2:0] n12445_o;
  wire [6:0] n12451_o;
  wire [3:0] n12453_o;
  wire n12455_o;
  wire n12456_o;
  wire n12457_o;
  wire n12459_o;
  wire n12460_o;
  wire n12462_o;
  wire n12465_o;
  wire n12467_o;
  wire [31:0] n12469_o;
  wire [5:0] n12470_o;
  wire n12472_o;
  wire [1:0] n12473_o;
  wire n12475_o;
  wire n12476_o;
  wire [4:0] n12477_o;
  wire n12479_o;
  wire n12480_o;
  wire n12482_o;
  wire n12483_o;
  wire n12485_o;
  wire n12486_o;
  wire n12488_o;
  wire n12489_o;
  wire n12491_o;
  wire n12493_o;
  wire n12495_o;
  wire [63:0] n12496_o;
  wire [5:0] n12497_o;
  wire [63:0] n12499_o;
  wire [31:0] n12501_o;
  wire [2:0] n12504_o;
  wire n12505_o;
  wire n12507_o;
  wire n12508_o;
  wire [1:0] n12509_o;
  wire [6:0] n12514_o;
  wire n12516_o;
  wire n12518_o;
  wire [798:0] n12519_o;
  wire [389:0] n12520_o;
  wire [63:0] n12523_o;
  wire [32:0] n12529_o;
  localparam [63:0] n12530_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire [4:0] n12532_o;
  wire [3:0] n12533_o;
  wire [15:0] n12535_o;
  wire [5:0] n12536_o;
  wire [63:0] n12537_o;
  wire [289:0] n12538_o;
  wire [309:0] n12539_o;
  reg [798:0] n12548_q;
  reg [255:0] n12549_q;
  wire [255:0] n12550_o;
  wire [258:0] n12553_o;
  wire [133:0] n12554_o;
  wire [227:0] n12555_o;
  wire [353:0] n12556_o;
  wire [66:0] n12557_o;
  wire [34:0] n12558_o;
  localparam [14:0] n12559_o = 15'bZ;
  wire n12561_data; // mem_rd
  wire n12562_o;
  wire n12563_o;
  wire n12564_o;
  wire n12565_o;
  wire n12566_o;
  wire n12567_o;
  wire n12568_o;
  wire n12569_o;
  wire n12570_o;
  wire n12571_o;
  wire n12572_o;
  wire n12573_o;
  wire n12574_o;
  wire n12575_o;
  wire n12576_o;
  wire n12577_o;
  wire n12578_o;
  wire n12579_o;
  wire n12580_o;
  wire n12581_o;
  wire n12582_o;
  wire n12583_o;
  wire n12584_o;
  wire n12585_o;
  wire n12586_o;
  wire n12587_o;
  wire n12588_o;
  wire n12589_o;
  wire n12590_o;
  wire n12591_o;
  wire n12592_o;
  wire n12593_o;
  wire [1:0] n12594_o;
  reg n12595_o;
  wire [1:0] n12596_o;
  reg n12597_o;
  wire [1:0] n12598_o;
  reg n12599_o;
  wire [1:0] n12600_o;
  reg n12601_o;
  wire [1:0] n12602_o;
  reg n12603_o;
  wire [1:0] n12604_o;
  reg n12605_o;
  wire [1:0] n12606_o;
  reg n12607_o;
  wire [1:0] n12608_o;
  reg n12609_o;
  wire [1:0] n12610_o;
  reg n12611_o;
  wire [1:0] n12612_o;
  reg n12613_o;
  wire n12614_o;
  wire n12615_o;
  wire n12616_o;
  wire n12617_o;
  wire n12618_o;
  wire n12619_o;
  wire n12620_o;
  wire n12621_o;
  wire n12622_o;
  wire n12623_o;
  wire n12624_o;
  wire n12625_o;
  wire n12626_o;
  wire n12627_o;
  wire n12628_o;
  wire n12629_o;
  wire n12630_o;
  wire n12631_o;
  wire n12632_o;
  wire n12633_o;
  wire n12634_o;
  wire n12635_o;
  wire n12636_o;
  wire n12637_o;
  wire n12638_o;
  wire n12639_o;
  wire n12640_o;
  wire n12641_o;
  wire n12642_o;
  wire n12643_o;
  wire n12644_o;
  wire n12645_o;
  wire n12646_o;
  wire n12647_o;
  wire [1:0] n12648_o;
  reg n12649_o;
  wire [1:0] n12650_o;
  reg n12651_o;
  wire [1:0] n12652_o;
  reg n12653_o;
  wire [1:0] n12654_o;
  reg n12655_o;
  wire [1:0] n12656_o;
  reg n12657_o;
  wire [1:0] n12658_o;
  reg n12659_o;
  wire [1:0] n12660_o;
  reg n12661_o;
  wire [1:0] n12662_o;
  reg n12663_o;
  wire [1:0] n12664_o;
  reg n12665_o;
  wire [1:0] n12666_o;
  reg n12667_o;
  wire n12668_o;
  wire n12669_o;
  wire n12670_o;
  wire n12671_o;
  wire n12672_o;
  wire n12673_o;
  wire n12674_o;
  wire n12675_o;
  wire n12676_o;
  wire n12677_o;
  wire n12678_o;
  wire n12679_o;
  wire n12680_o;
  wire n12681_o;
  wire n12682_o;
  wire n12683_o;
  wire n12684_o;
  wire n12685_o;
  wire n12686_o;
  wire n12687_o;
  wire n12688_o;
  wire n12689_o;
  wire n12690_o;
  wire n12691_o;
  wire n12692_o;
  wire n12693_o;
  wire n12694_o;
  wire n12695_o;
  wire n12696_o;
  wire n12697_o;
  wire n12698_o;
  wire n12699_o;
  wire n12700_o;
  wire n12701_o;
  wire [1:0] n12702_o;
  reg n12703_o;
  wire [1:0] n12704_o;
  reg n12705_o;
  wire [1:0] n12706_o;
  reg n12707_o;
  wire [1:0] n12708_o;
  reg n12709_o;
  wire [1:0] n12710_o;
  reg n12711_o;
  wire [1:0] n12712_o;
  reg n12713_o;
  wire [1:0] n12714_o;
  reg n12715_o;
  wire [1:0] n12716_o;
  reg n12717_o;
  wire [1:0] n12718_o;
  reg n12719_o;
  wire [1:0] n12720_o;
  reg n12721_o;
  wire n12722_o;
  wire n12723_o;
  wire [3:0] n12724_o;
  wire [3:0] n12725_o;
  wire [3:0] n12726_o;
  wire [3:0] n12727_o;
  wire [3:0] n12728_o;
  wire [3:0] n12729_o;
  wire [3:0] n12730_o;
  wire [3:0] n12731_o;
  wire [1:0] n12732_o;
  reg [3:0] n12733_o;
  wire [1:0] n12734_o;
  reg [3:0] n12735_o;
  wire n12736_o;
  wire [3:0] n12737_o;
  wire n12738_o;
  wire n12739_o;
  wire n12740_o;
  wire n12741_o;
  wire n12742_o;
  wire n12743_o;
  wire n12744_o;
  wire n12745_o;
  wire n12746_o;
  wire n12747_o;
  wire n12748_o;
  wire n12749_o;
  wire n12750_o;
  wire n12751_o;
  wire n12752_o;
  wire n12753_o;
  wire n12754_o;
  wire n12755_o;
  wire n12756_o;
  wire n12757_o;
  wire n12758_o;
  wire n12759_o;
  wire n12760_o;
  wire n12761_o;
  wire n12762_o;
  wire n12763_o;
  wire n12764_o;
  wire n12765_o;
  wire n12766_o;
  wire n12767_o;
  wire n12768_o;
  wire n12769_o;
  wire [1:0] n12770_o;
  reg n12771_o;
  wire [1:0] n12772_o;
  reg n12773_o;
  wire [1:0] n12774_o;
  reg n12775_o;
  wire [1:0] n12776_o;
  reg n12777_o;
  wire [1:0] n12778_o;
  reg n12779_o;
  wire [1:0] n12780_o;
  reg n12781_o;
  wire [1:0] n12782_o;
  reg n12783_o;
  wire [1:0] n12784_o;
  reg n12785_o;
  wire [1:0] n12786_o;
  reg n12787_o;
  wire [1:0] n12788_o;
  reg n12789_o;
  wire n12790_o;
  wire n12791_o;
  wire n12792_o;
  wire n12793_o;
  wire n12794_o;
  wire n12795_o;
  wire n12796_o;
  wire n12797_o;
  wire n12798_o;
  wire n12799_o;
  wire n12800_o;
  wire n12801_o;
  wire n12802_o;
  wire n12803_o;
  wire n12804_o;
  wire n12805_o;
  wire n12806_o;
  wire n12807_o;
  wire n12808_o;
  wire n12809_o;
  wire n12810_o;
  wire n12811_o;
  wire n12812_o;
  wire n12813_o;
  wire n12814_o;
  wire n12815_o;
  wire n12816_o;
  wire n12817_o;
  wire n12818_o;
  wire n12819_o;
  wire n12820_o;
  wire n12821_o;
  wire n12822_o;
  wire n12823_o;
  wire [1:0] n12824_o;
  reg n12825_o;
  wire [1:0] n12826_o;
  reg n12827_o;
  wire [1:0] n12828_o;
  reg n12829_o;
  wire [1:0] n12830_o;
  reg n12831_o;
  wire [1:0] n12832_o;
  reg n12833_o;
  wire [1:0] n12834_o;
  reg n12835_o;
  wire [1:0] n12836_o;
  reg n12837_o;
  wire [1:0] n12838_o;
  reg n12839_o;
  wire [1:0] n12840_o;
  reg n12841_o;
  wire [1:0] n12842_o;
  reg n12843_o;
  wire n12844_o;
  wire n12845_o;
  wire n12846_o;
  wire n12847_o;
  wire n12848_o;
  wire n12849_o;
  wire n12850_o;
  wire n12851_o;
  wire n12852_o;
  wire n12853_o;
  wire n12854_o;
  wire n12855_o;
  wire n12856_o;
  wire n12857_o;
  wire n12858_o;
  wire n12859_o;
  wire n12860_o;
  wire n12861_o;
  wire n12862_o;
  wire n12863_o;
  wire n12864_o;
  wire n12865_o;
  wire n12866_o;
  wire n12867_o;
  wire n12868_o;
  wire n12869_o;
  wire n12870_o;
  wire n12871_o;
  wire n12872_o;
  wire n12873_o;
  wire n12874_o;
  wire n12875_o;
  wire n12876_o;
  wire n12877_o;
  wire [1:0] n12878_o;
  reg n12879_o;
  wire [1:0] n12880_o;
  reg n12881_o;
  wire [1:0] n12882_o;
  reg n12883_o;
  wire [1:0] n12884_o;
  reg n12885_o;
  wire [1:0] n12886_o;
  reg n12887_o;
  wire [1:0] n12888_o;
  reg n12889_o;
  wire [1:0] n12890_o;
  reg n12891_o;
  wire [1:0] n12892_o;
  reg n12893_o;
  wire [1:0] n12894_o;
  reg n12895_o;
  wire [1:0] n12896_o;
  reg n12897_o;
  wire n12898_o;
  wire n12899_o;
  wire [3:0] n12900_o;
  wire [3:0] n12901_o;
  wire [3:0] n12902_o;
  wire [3:0] n12903_o;
  wire [3:0] n12904_o;
  wire [3:0] n12905_o;
  wire [3:0] n12906_o;
  wire [3:0] n12907_o;
  wire [1:0] n12908_o;
  reg [3:0] n12909_o;
  wire [1:0] n12910_o;
  reg [3:0] n12911_o;
  wire n12912_o;
  wire [3:0] n12913_o;
  wire n12914_o;
  wire n12915_o;
  wire n12916_o;
  wire n12917_o;
  wire n12918_o;
  wire n12919_o;
  wire n12920_o;
  wire n12921_o;
  wire n12922_o;
  wire n12923_o;
  wire n12924_o;
  wire n12925_o;
  wire n12926_o;
  wire n12927_o;
  wire n12928_o;
  wire n12929_o;
  wire n12930_o;
  wire n12931_o;
  wire n12932_o;
  wire n12933_o;
  wire n12934_o;
  wire n12935_o;
  wire n12936_o;
  wire n12937_o;
  wire n12938_o;
  wire n12939_o;
  wire n12940_o;
  wire n12941_o;
  wire n12942_o;
  wire n12943_o;
  wire n12944_o;
  wire n12945_o;
  wire [1:0] n12946_o;
  reg n12947_o;
  wire [1:0] n12948_o;
  reg n12949_o;
  wire [1:0] n12950_o;
  reg n12951_o;
  wire [1:0] n12952_o;
  reg n12953_o;
  wire [1:0] n12954_o;
  reg n12955_o;
  wire [1:0] n12956_o;
  reg n12957_o;
  wire [1:0] n12958_o;
  reg n12959_o;
  wire [1:0] n12960_o;
  reg n12961_o;
  wire [1:0] n12962_o;
  reg n12963_o;
  wire [1:0] n12964_o;
  reg n12965_o;
  wire n12966_o;
  wire n12967_o;
  assign busy_out = n9336_o;
  assign l_out_valid = n9143_o;
  assign l_out_op = n9144_o;
  assign l_out_nia = n9145_o;
  assign l_out_insn = n9146_o;
  assign l_out_instr_tag = n9147_o;
  assign l_out_addr1 = n9148_o;
  assign l_out_addr2 = n9149_o;
  assign l_out_data = n9150_o;
  assign l_out_write_reg = n9151_o;
  assign l_out_length = n9152_o;
  assign l_out_ci = n9153_o;
  assign l_out_byte_reverse = n9154_o;
  assign l_out_sign_extend = n9155_o;
  assign l_out_update = n9156_o;
  assign l_out_xerc = n9157_o;
  assign l_out_reserve = n9158_o;
  assign l_out_rc = n9159_o;
  assign l_out_virt_mode = n9160_o;
  assign l_out_priv_mode = n9161_o;
  assign l_out_mode_32bit = n9162_o;
  assign l_out_is_32bit = n9163_o;
  assign l_out_repeat = n9164_o;
  assign l_out_second = n9165_o;
  assign l_out_msr = n9166_o;
  assign fp_out_valid = n9168_o;
  assign fp_out_op = n9169_o;
  assign fp_out_nia = n9170_o;
  assign fp_out_itag = n9171_o;
  assign fp_out_insn = n9172_o;
  assign fp_out_single = n9173_o;
  assign fp_out_fe_mode = n9174_o;
  assign fp_out_fra = n9175_o;
  assign fp_out_frb = n9176_o;
  assign fp_out_frc = n9177_o;
  assign fp_out_frt = n9178_o;
  assign fp_out_rc = n9179_o;
  assign fp_out_out_cr = n9180_o;
  assign e_out_valid = n9182_o;
  assign e_out_instr_tag = n9183_o;
  assign e_out_rc = n9184_o;
  assign e_out_mode_32bit = n9185_o;
  assign e_out_write_enable = n9186_o;
  assign e_out_write_reg = n9187_o;
  assign e_out_write_data = n9188_o;
  assign e_out_write_cr_enable = n9189_o;
  assign e_out_write_cr_mask = n9190_o;
  assign e_out_write_cr_data = n9191_o;
  assign e_out_write_xerc_enable = n9192_o;
  assign e_out_xerc = n9193_o;
  assign e_out_interrupt = n9194_o;
  assign e_out_intr_vec = n9195_o;
  assign e_out_redirect = n9196_o;
  assign e_out_redir_mode = n9197_o;
  assign e_out_last_nia = n9198_o;
  assign e_out_br_offset = n9199_o;
  assign e_out_br_last = n9200_o;
  assign e_out_br_taken = n9201_o;
  assign e_out_abs_br = n9202_o;
  assign e_out_srr1 = n9203_o;
  assign e_out_msr = n9204_o;
  assign bypass_data_tag = n9206_o;
  assign bypass_data_data = n9207_o;
  assign bypass_cr_data_tag = n9209_o;
  assign bypass_cr_data_data = n9210_o;
  assign dbg_msr_out = n9273_o;
  assign icache_inval = n11992_o;
  assign terminate_out = n9342_o;
  assign log_out = n12559_o;
  assign log_rd_addr = n9274_o;
  /* common.vhdl:112:14  */
  assign n9139_o = {e_in_second, e_in_repeat, e_in_sub_select, e_in_result_sel, e_in_br_pred, e_in_reserve, e_in_update, e_in_sign_extend, e_in_byte_reverse, e_in_data_len, e_in_insn, e_in_is_signed, e_in_is_32bit, e_in_output_xer, e_in_output_cr, e_in_input_cr, e_in_output_carry, e_in_input_carry, e_in_invert_out, e_in_addm1, e_in_invert_a, e_in_oe, e_in_rc, e_in_br_abs, e_in_lr, e_in_xerc, e_in_cr, e_in_read_data3, e_in_read_data2, e_in_read_data1, e_in_read_reg2, e_in_read_reg1, e_in_write_reg_enable, e_in_write_reg, e_in_instr_tag, e_in_nia, e_in_insn_type, e_in_fac, e_in_unit, e_in_valid};
  /* cr_file.vhdl:78:17  */
  assign n9140_o = {l_in_interrupt, l_in_in_progress, l_in_busy};
  /* cr_file.vhdl:75:5  */
  assign n9141_o = {fp_in_exception, fp_in_busy};
  /* cr_file.vhdl:62:9  */
  assign n9143_o = n12520_o[0];
  /* cr_file.vhdl:62:9  */
  assign n9144_o = n12520_o[6:1];
  /* cr_file.vhdl:60:5  */
  assign n9145_o = n12520_o[70:7];
  /* insn_helpers.vhdl:5:14  */
  assign n9146_o = n12520_o[102:71];
  /* common.vhdl:110:14  */
  assign n9147_o = n12520_o[105:103];
  /* cr_file.vhdl:42:13  */
  assign n9148_o = n12520_o[169:106];
  /* insn_helpers.vhdl:9:14  */
  assign n9149_o = n12520_o[233:170];
  /* cr_file.vhdl:42:13  */
  assign n9150_o = n12520_o[297:234];
  assign n9151_o = n12520_o[304:298];
  /* cr_file.vhdl:42:13  */
  assign n9152_o = n12520_o[308:305];
  /* common.vhdl:113:14  */
  assign n9153_o = n12520_o[309];
  /* cr_file.vhdl:42:13  */
  assign n9154_o = n12520_o[310];
  /* common.vhdl:113:14  */
  assign n9155_o = n12520_o[311];
  assign n9156_o = n12520_o[312];
  /* cr_file.vhdl:42:13  */
  assign n9157_o = n12520_o[317:313];
  assign n9158_o = n12520_o[318];
  /* cr_file.vhdl:42:13  */
  assign n9159_o = n12520_o[319];
  /* common.vhdl:113:14  */
  assign n9160_o = n12520_o[320];
  /* decode2.vhdl:172:14  */
  assign n9161_o = n12520_o[321];
  /* cr_file.vhdl:42:13  */
  assign n9162_o = n12520_o[322];
  /* insn_helpers.vhdl:6:14  */
  assign n9163_o = n12520_o[323];
  /* cr_file.vhdl:42:13  */
  assign n9164_o = n12520_o[324];
  /* common.vhdl:110:14  */
  assign n9165_o = n12520_o[325];
  /* common.vhdl:110:14  */
  assign n9166_o = n12520_o[389:326];
  /* insn_helpers.vhdl:7:14  */
  assign n9168_o = n12539_o[0];
  /* cr_file.vhdl:42:13  */
  assign n9169_o = n12539_o[6:1];
  assign n9170_o = n12539_o[70:7];
  /* insn_helpers.vhdl:41:14  */
  assign n9171_o = n12539_o[73:71];
  /* cr_file.vhdl:42:13  */
  assign n9172_o = n12539_o[105:74];
  /* common.vhdl:113:14  */
  assign n9173_o = n12539_o[106];
  /* cr_file.vhdl:42:13  */
  assign n9174_o = n12539_o[108:107];
  /* common.vhdl:113:14  */
  assign n9175_o = n12539_o[172:109];
  assign n9176_o = n12539_o[236:173];
  /* cr_file.vhdl:42:13  */
  assign n9177_o = n12539_o[300:237];
  assign n9178_o = n12539_o[307:301];
  /* cr_file.vhdl:42:13  */
  assign n9179_o = n12539_o[308];
  /* insn_helpers.vhdl:17:14  */
  assign n9180_o = n12539_o[309];
  /* cr_file.vhdl:42:13  */
  assign n9182_o = n12556_o[0];
  assign n9183_o = n12556_o[3:1];
  /* cr_file.vhdl:42:13  */
  assign n9184_o = n12556_o[4];
  assign n9185_o = n12556_o[5];
  /* cr_file.vhdl:35:5  */
  assign n9186_o = n12556_o[6];
  /* cr_file.vhdl:37:18  */
  assign n9187_o = n12556_o[13:7];
  assign n9188_o = n12556_o[77:14];
  /* cr_file.vhdl:36:22  */
  assign n9189_o = n12556_o[78];
  /* decode2.vhdl:199:14  */
  assign n9190_o = n12556_o[86:79];
  /* cr_file.vhdl:36:18  */
  assign n9191_o = n12556_o[118:87];
  /* asic/register_file.vhdl:76:12  */
  assign n9192_o = n12556_o[119];
  /* insn_helpers.vhdl:34:14  */
  assign n9193_o = n12556_o[124:120];
  /* insn_helpers.vhdl:34:14  */
  assign n9194_o = n12556_o[125];
  assign n9195_o = n12556_o[137:126];
  /* insn_helpers.vhdl:34:14  */
  assign n9196_o = n12556_o[138];
  /* insn_helpers.vhdl:33:14  */
  assign n9197_o = n12556_o[142:139];
  /* insn_helpers.vhdl:33:14  */
  assign n9198_o = n12556_o[206:143];
  assign n9199_o = n12556_o[270:207];
  /* insn_helpers.vhdl:33:14  */
  assign n9200_o = n12556_o[271];
  /* insn_helpers.vhdl:21:14  */
  assign n9201_o = n12556_o[272];
  /* insn_helpers.vhdl:21:14  */
  assign n9202_o = n12556_o[273];
  assign n9203_o = n12556_o[289:274];
  /* insn_helpers.vhdl:21:14  */
  assign n9204_o = n12556_o[353:290];
  /* insn_helpers.vhdl:16:14  */
  assign n9206_o = n12557_o[2:0];
  assign n9207_o = n12557_o[66:3];
  /* insn_helpers.vhdl:10:14  */
  assign n9209_o = n12558_o[2:0];
  /* insn_helpers.vhdl:10:14  */
  assign n9210_o = n12558_o[34:3];
  /* insn_helpers.vhdl:10:14  */
  assign n9214_o = {wb_events_fp_complete, wb_events_instr_complete};
  assign n9215_o = {ls_events_itlb_miss, ls_events_store_complete, ls_events_load_complete};
  /* insn_helpers.vhdl:10:14  */
  assign n9216_o = {dc_events_dtlb_miss_resolved, dc_events_dtlb_miss, dc_events_dcache_refill, dc_events_store_miss, dc_events_load_miss};
  /* insn_helpers.vhdl:10:14  */
  assign n9217_o = {ic_events_itlb_miss_resolved, ic_events_icache_miss};
  /* execute1.vhdl:94:12  */
  assign r = n12548_q; // (signal)
  /* execute1.vhdl:94:15  */
  assign rin = n12519_o; // (signal)
  /* execute1.vhdl:96:12  */
  assign a_in = n9275_o; // (signal)
  /* execute1.vhdl:96:18  */
  assign b_in = n9276_o; // (signal)
  /* execute1.vhdl:96:24  */
  assign c_in = n9277_o; // (signal)
  /* execute1.vhdl:97:12  */
  assign cr_in = n9278_o; // (signal)
  /* execute1.vhdl:98:12  */
  assign xerc_in = n9319_o; // (signal)
  /* execute1.vhdl:101:12  */
  assign valid_in = n9341_o; // (signal)
  /* execute1.vhdl:102:12  */
  always @*
    ctrl = n12549_q; // (isignal)
  initial
    ctrl = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* execute1.vhdl:103:12  */
  always @*
    ctrl_tmp = n12550_o; // (isignal)
  initial
    ctrl_tmp = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* execute1.vhdl:104:12  */
  assign right_shift = n10772_o; // (signal)
  /* execute1.vhdl:104:25  */
  assign rot_clear_left = n10782_o; // (signal)
  /* execute1.vhdl:104:41  */
  assign rot_clear_right = n10792_o; // (signal)
  /* execute1.vhdl:105:12  */
  assign rot_sign_ext = n10798_o; // (signal)
  /* execute1.vhdl:106:12  */
  assign rotator_result = rotator_0_result; // (signal)
  /* execute1.vhdl:107:12  */
  assign rotator_carry = rotator_0_carry_out; // (signal)
  /* execute1.vhdl:108:12  */
  assign logical_result = logical_0_result; // (signal)
  /* execute1.vhdl:109:12  */
  assign do_popcnt = n10804_o; // (signal)
  /* execute1.vhdl:110:12  */
  assign countbits_result = countbits_0_result; // (signal)
  /* execute1.vhdl:111:12  */
  assign alu_result = n9363_o; // (signal)
  /* execute1.vhdl:112:12  */
  assign adder_result = n9459_o; // (signal)
  /* execute1.vhdl:113:12  */
  assign misc_result = n10097_o; // (signal)
  /* execute1.vhdl:114:12  */
  assign muldiv_result = n9670_o; // (signal)
  /* execute1.vhdl:115:12  */
  assign spr_result = n11998_o; // (signal)
  /* execute1.vhdl:118:12  */
  assign next_nia = n10767_o; // (signal)
  /* execute1.vhdl:119:12  */
  assign current = n9345_o; // (signal)
  /* execute1.vhdl:121:12  */
  assign carry_32 = n9464_o; // (signal)
  /* execute1.vhdl:122:12  */
  assign carry_64 = n9465_o; // (signal)
  /* execute1.vhdl:123:12  */
  assign overflow_32 = n9477_o; // (signal)
  /* execute1.vhdl:124:12  */
  assign overflow_64 = n9489_o; // (signal)
  /* execute1.vhdl:126:12  */
  assign trapval = n10212_o; // (signal)
  /* execute1.vhdl:128:12  */
  assign write_cr_mask = n10680_o; // (signal)
  /* execute1.vhdl:129:12  */
  assign write_cr_data = n10681_o; // (signal)
  /* execute1.vhdl:132:12  */
  assign x_to_multiply = n12553_o; // (signal)
  /* execute1.vhdl:133:12  */
  assign multiply_to_x = n9244_o; // (signal)
  /* execute1.vhdl:136:12  */
  assign x_to_divider = n12554_o; // (signal)
  /* execute1.vhdl:137:12  */
  assign divider_to_x = n9254_o; // (signal)
  /* execute1.vhdl:140:12  */
  assign random_raw = random_0_raw; // (signal)
  /* execute1.vhdl:141:12  */
  assign random_cond = random_0_data; // (signal)
  /* execute1.vhdl:142:12  */
  assign random_err = random_0_err; // (signal)
  /* execute1.vhdl:145:12  */
  assign x_to_pmu = n12555_o; // (signal)
  /* execute1.vhdl:146:12  */
  assign pmu_to_x = n9271_o; // (signal)
  /* execute1.vhdl:261:5  */
  rotator rotator_0 (
    .rs(c_in),
    .ra(a_in),
    .shift(n9223_o),
    .insn(n9224_o),
    .is_32bit(n9225_o),
    .right_shift(right_shift),
    .arith(n9226_o),
    .clear_left(rot_clear_left),
    .clear_right(rot_clear_right),
    .sign_ext_rs(rot_sign_ext),
    .result(rotator_0_result),
    .carry_out(rotator_0_carry_out));
  /* execute1.vhdl:265:26  */
  assign n9223_o = b_in[6:0];
  /* execute1.vhdl:266:26  */
  assign n9224_o = n9139_o[374:343];
  /* execute1.vhdl:267:30  */
  assign n9225_o = n9139_o[341];
  /* execute1.vhdl:269:27  */
  assign n9226_o = n9139_o[342];
  /* execute1.vhdl:277:5  */
  logical logical_0 (
    .rs(c_in),
    .rb(b_in),
    .op(n9229_o),
    .invert_in(n9230_o),
    .invert_out(n9231_o),
    .datalen(n9233_o),
    .result(logical_0_result));
  /* execute1.vhdl:281:24  */
  assign n9229_o = n9139_o[9:4];
  /* execute1.vhdl:282:31  */
  assign n9230_o = n9139_o[332];
  /* execute1.vhdl:283:32  */
  assign n9231_o = n9139_o[334];
  /* execute1.vhdl:285:29  */
  assign n9233_o = n9139_o[378:375];
  /* execute1.vhdl:288:5  */
  bit_counter countbits_0 (
    .clk(clk),
    .rs(c_in),
    .count_right(n9234_o),
    .do_popcnt(do_popcnt),
    .is_32bit(n9235_o),
    .datalen(n9236_o),
    .result(countbits_0_result));
  /* execute1.vhdl:292:37  */
  assign n9234_o = n9139_o[353];
  /* execute1.vhdl:293:30  */
  assign n9235_o = n9139_o[341];
  /* execute1.vhdl:295:29  */
  assign n9236_o = n9139_o[378:375];
  /* execute1.vhdl:299:5  */
  multiply_2 multiply_0 (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(clk),
    .m_in_valid(n9238_o),
    .m_in_data1(n9239_o),
    .m_in_data2(n9240_o),
    .m_in_addend(n9241_o),
    .m_in_is_32bit(n9242_o),
    .m_in_not_result(n9243_o),
    .m_out_valid(multiply_0_m_out_valid),
    .m_out_result(multiply_0_m_out_result),
    .m_out_overflow(multiply_0_m_out_overflow));
  assign n9238_o = x_to_multiply[0];
  /* decode2.vhdl:372:18  */
  assign n9239_o = x_to_multiply[64:1];
  assign n9240_o = x_to_multiply[128:65];
  /* decode2.vhdl:371:18  */
  assign n9241_o = x_to_multiply[256:129];
  assign n9242_o = x_to_multiply[257];
  /* decode2.vhdl:370:18  */
  assign n9243_o = x_to_multiply[258];
  assign n9244_o = {multiply_0_m_out_overflow, multiply_0_m_out_result, multiply_0_m_out_valid};
  /* execute1.vhdl:306:5  */
  divider divider_0 (
    .clk(clk),
    .rst(rst),
    .d_in_valid(n9246_o),
    .d_in_dividend(n9247_o),
    .d_in_divisor(n9248_o),
    .d_in_is_signed(n9249_o),
    .d_in_is_32bit(n9250_o),
    .d_in_is_extended(n9251_o),
    .d_in_is_modulus(n9252_o),
    .d_in_neg_result(n9253_o),
    .d_out_valid(divider_0_d_out_valid),
    .d_out_write_reg_data(divider_0_d_out_write_reg_data),
    .d_out_overflow(divider_0_d_out_overflow));
  /* decode2.vhdl:368:18  */
  assign n9246_o = x_to_divider[0];
  assign n9247_o = x_to_divider[64:1];
  /* decode2.vhdl:367:18  */
  assign n9248_o = x_to_divider[128:65];
  assign n9249_o = x_to_divider[129];
  /* decode2.vhdl:366:18  */
  assign n9250_o = x_to_divider[130];
  assign n9251_o = x_to_divider[131];
  /* decode2.vhdl:365:18  */
  assign n9252_o = x_to_divider[132];
  assign n9253_o = x_to_divider[133];
  assign n9254_o = {divider_0_d_out_overflow, divider_0_d_out_write_reg_data, divider_0_d_out_valid};
  /* execute1.vhdl:314:5  */
  random random_0 (
    .clk(clk),
    .data(random_0_data),
    .raw(random_0_raw),
    .err(random_0_err));
  /* execute1.vhdl:322:5  */
  pmu pmu_0 (
    .clk(clk),
    .rst(rst),
    .p_in_mfspr(n9259_o),
    .p_in_mtspr(n9260_o),
    .p_in_spr_num(n9261_o),
    .p_in_spr_val(n9262_o),
    .p_in_tbbits(n9263_o),
    .p_in_pmm_msr(n9264_o),
    .p_in_pr_msr(n9265_o),
    .p_in_run(n9266_o),
    .p_in_nia(n9267_o),
    .p_in_addr(n9268_o),
    .p_in_addr_v(n9269_o),
    .p_in_occur(n9270_o),
    .p_out_spr_val(pmu_0_p_out_spr_val),
    .p_out_intr(pmu_0_p_out_intr));
  assign n9259_o = x_to_pmu[0];
  assign n9260_o = x_to_pmu[1];
  assign n9261_o = x_to_pmu[6:2];
  assign n9262_o = x_to_pmu[70:7];
  assign n9263_o = x_to_pmu[74:71];
  assign n9264_o = x_to_pmu[75];
  assign n9265_o = x_to_pmu[76];
  assign n9266_o = x_to_pmu[77];
  assign n9267_o = x_to_pmu[141:78];
  assign n9268_o = x_to_pmu[205:142];
  assign n9269_o = x_to_pmu[206];
  assign n9270_o = x_to_pmu[227:207];
  assign n9271_o = {pmu_0_p_out_intr, pmu_0_p_out_spr_val};
  /* execute1.vhdl:341:25  */
  assign n9273_o = ctrl[191:128];
  /* execute1.vhdl:342:22  */
  assign n9274_o = r[798:767];
  /* execute1.vhdl:344:18  */
  assign n9275_o = n9139_o[162:99];
  /* execute1.vhdl:345:18  */
  assign n9276_o = n9139_o[226:163];
  /* execute1.vhdl:346:18  */
  assign n9277_o = n9139_o[290:227];
  /* execute1.vhdl:347:19  */
  assign n9278_o = n9139_o[322:291];
  /* execute1.vhdl:349:52  */
  assign n9279_o = n9214_o[0];
  /* execute1.vhdl:350:49  */
  assign n9280_o = n9214_o[1];
  /* execute1.vhdl:351:49  */
  assign n9281_o = n9215_o[0];
  /* execute1.vhdl:352:49  */
  assign n9282_o = n9215_o[1];
  /* execute1.vhdl:353:47  */
  assign n9283_o = n9215_o[2];
  /* execute1.vhdl:354:50  */
  assign n9284_o = n9216_o[0];
  /* execute1.vhdl:355:57  */
  assign n9285_o = n9216_o[2];
  /* execute1.vhdl:356:51  */
  assign n9286_o = n9216_o[1];
  /* execute1.vhdl:357:47  */
  assign n9287_o = n9216_o[3];
  /* execute1.vhdl:358:56  */
  assign n9288_o = n9216_o[4];
  /* execute1.vhdl:359:49  */
  assign n9289_o = n9217_o[0];
  /* execute1.vhdl:360:56  */
  assign n9290_o = n9217_o[1];
  /* execute1.vhdl:361:44  */
  assign n9291_o = r[762];
  /* execute1.vhdl:362:38  */
  assign n9292_o = r[763];
  /* execute1.vhdl:363:43  */
  assign n9293_o = r[764];
  /* execute1.vhdl:364:47  */
  assign n9294_o = r[765];
  /* execute1.vhdl:365:43  */
  assign n9295_o = r[766];
  assign n9300_o = {1'b0, 1'b0, n9288_o, n9287_o};
  assign n9301_o = {n9286_o, n9285_o, n9284_o, 1'b0};
  assign n9302_o = {n9289_o, n9290_o, n9283_o, 1'b0};
  assign n9303_o = {n9295_o, n9294_o, n9282_o, n9281_o};
  assign n9304_o = {n9280_o, n9279_o, n9293_o, n9292_o};
  assign n9305_o = {n9300_o, n9301_o, n9302_o, n9303_o};
  assign n9306_o = {n9304_o, n9291_o};
  assign n9307_o = {n9305_o, n9306_o};
  /* execute1.vhdl:367:29  */
  assign n9308_o = current[73:10];
  /* execute1.vhdl:370:34  */
  assign n9311_o = n9139_o[363:359];
  /* execute1.vhdl:379:18  */
  assign n9313_o = r[353:0];
  /* execute1.vhdl:379:20  */
  assign n9314_o = n9313_o[124:120];
  /* execute1.vhdl:379:32  */
  assign n9315_o = r[353:0];
  /* execute1.vhdl:379:34  */
  assign n9316_o = n9315_o[119];
  /* execute1.vhdl:379:63  */
  assign n9317_o = r[746];
  /* execute1.vhdl:379:58  */
  assign n9318_o = n9316_o | n9317_o;
  /* execute1.vhdl:379:25  */
  assign n9319_o = n9318_o ? n9314_o : n9320_o;
  /* execute1.vhdl:379:84  */
  assign n9320_o = n9139_o[327:323];
  /* execute1.vhdl:381:15  */
  assign n9321_o = n9139_o[2:1];
  /* execute1.vhdl:382:14  */
  assign n9322_o = n9140_o[0];
  /* execute1.vhdl:382:24  */
  assign n9323_o = r[746];
  /* execute1.vhdl:382:19  */
  assign n9324_o = n9322_o | n9323_o;
  /* execute1.vhdl:382:38  */
  assign n9325_o = n9141_o[0];
  /* execute1.vhdl:382:29  */
  assign n9326_o = n9324_o | n9325_o;
  /* execute1.vhdl:382:43  */
  assign n9328_o = n9321_o == 2'b10;
  /* execute1.vhdl:383:14  */
  assign n9329_o = n9140_o[0];
  /* execute1.vhdl:383:27  */
  assign n9330_o = n9140_o[1];
  /* execute1.vhdl:383:19  */
  assign n9331_o = n9329_o | n9330_o;
  /* execute1.vhdl:383:44  */
  assign n9332_o = r[746];
  /* execute1.vhdl:383:39  */
  assign n9333_o = n9331_o | n9332_o;
  /* execute1.vhdl:383:58  */
  assign n9334_o = n9141_o[0];
  /* execute1.vhdl:383:49  */
  assign n9335_o = n9333_o | n9334_o;
  /* execute1.vhdl:381:5  */
  always @*
    case (n9328_o)
      1'b1: n9336_o = n9326_o;
      default: n9336_o = n9335_o;
    endcase
  /* execute1.vhdl:385:22  */
  assign n9337_o = n9139_o[0];
  /* execute1.vhdl:385:32  */
  assign n9338_o = ~n9336_o;
  /* execute1.vhdl:385:28  */
  assign n9339_o = n9337_o & n9338_o;
  /* execute1.vhdl:385:49  */
  assign n9340_o = ~flush_in;
  /* execute1.vhdl:385:45  */
  assign n9341_o = n9339_o & n9340_o;
  /* execute1.vhdl:387:24  */
  assign n9342_o = r[747];
  /* execute1.vhdl:389:28  */
  assign n9343_o = r[746];
  /* execute1.vhdl:389:33  */
  assign n9344_o = ~n9343_o;
  /* execute1.vhdl:389:21  */
  assign n9345_o = n9344_o ? n9139_o : n9346_o;
  /* execute1.vhdl:389:46  */
  assign n9346_o = r[745:354];
  /* execute1.vhdl:392:18  */
  assign n9347_o = current[386:384];
  /* execute1.vhdl:393:28  */
  assign n9349_o = n9347_o == 3'b000;
  /* execute1.vhdl:394:28  */
  assign n9351_o = n9347_o == 3'b001;
  /* execute1.vhdl:395:28  */
  assign n9353_o = n9347_o == 3'b010;
  /* execute1.vhdl:396:28  */
  assign n9355_o = n9347_o == 3'b011;
  /* execute1.vhdl:397:28  */
  assign n9357_o = n9347_o == 3'b100;
  /* execute1.vhdl:398:28  */
  assign n9359_o = n9347_o == 3'b101;
  /* execute1.vhdl:399:28  */
  assign n9361_o = n9347_o == 3'b110;
  assign n9362_o = {n9361_o, n9359_o, n9357_o, n9355_o, n9353_o, n9351_o, n9349_o};
  /* execute1.vhdl:392:5  */
  always @*
    case (n9362_o)
      7'b1000000: n9363_o = next_nia;
      7'b0100000: n9363_o = spr_result;
      7'b0010000: n9363_o = countbits_result;
      7'b0001000: n9363_o = muldiv_result;
      7'b0000100: n9363_o = rotator_result;
      7'b0000010: n9363_o = logical_result;
      7'b0000001: n9363_o = adder_result;
      default: n9363_o = misc_result;
    endcase
  /* execute1.vhdl:405:13  */
  assign n9370_o = rst ? 799'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : rin;
  assign n9371_o = {64'b1000000000000000000000000000000000000000000000000000000000000001, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000};
  assign n9372_o = ctrl_tmp[191:0];
  /* execute1.vhdl:405:13  */
  assign n9373_o = rst ? n9371_o : n9372_o;
  assign n9374_o = ctrl_tmp[255:192];
  assign n9375_o = ctrl[255:192];
  /* execute1.vhdl:405:13  */
  assign n9376_o = rst ? n9375_o : n9374_o;
  assign n9378_o = {n9376_o, n9373_o};
  /* execute1.vhdl:455:17  */
  assign n9420_o = n9139_o[332];
  /* execute1.vhdl:455:26  */
  assign n9421_o = ~n9420_o;
  /* execute1.vhdl:458:22  */
  assign n9422_o = ~a_in;
  /* execute1.vhdl:455:9  */
  assign n9423_o = n9421_o ? a_in : n9422_o;
  /* execute1.vhdl:460:17  */
  assign n9424_o = n9139_o[333];
  /* execute1.vhdl:460:23  */
  assign n9425_o = ~n9424_o;
  /* execute1.vhdl:460:9  */
  assign n9427_o = n9425_o ? b_in : 64'b1111111111111111111111111111111111111111111111111111111111111111;
  /* execute1.vhdl:466:60  */
  assign n9430_o = n9139_o[336:335];
  /* execute1.vhdl:204:9  */
  assign n9437_o = n9430_o == 2'b00;
  /* execute1.vhdl:207:25  */
  assign n9438_o = xerc_in[0];
  /* execute1.vhdl:206:9  */
  assign n9440_o = n9430_o == 2'b01;
  /* execute1.vhdl:209:25  */
  assign n9441_o = xerc_in[2];
  /* execute1.vhdl:208:9  */
  assign n9443_o = n9430_o == 2'b10;
  /* execute1.vhdl:210:9  */
  assign n9446_o = n9430_o == 2'b11;
  assign n9447_o = {n9446_o, n9443_o, n9440_o, n9437_o};
  /* execute1.vhdl:203:9  */
  always @*
    case (n9447_o)
      4'b1000: n9449_o = 1'b1;
      4'b0100: n9449_o = n9441_o;
      4'b0010: n9449_o = n9438_o;
      4'b0001: n9449_o = 1'b0;
      default: n9449_o = 1'bX;
    endcase
  /* ppc_fx_insns.vhdl:114:41  */
  assign n9454_o = {1'b0, n9423_o};  //  uext
  /* ppc_fx_insns.vhdl:114:68  */
  assign n9455_o = {1'b0, n9427_o};  //  uext
  /* ppc_fx_insns.vhdl:114:66  */
  assign n9456_o = n9454_o + n9455_o;
  /* ppc_fx_insns.vhdl:114:93  */
  assign n9457_o = {64'b0, n9449_o};  //  uext
  /* ppc_fx_insns.vhdl:114:93  */
  assign n9458_o = n9456_o + n9457_o;
  /* execute1.vhdl:467:39  */
  assign n9459_o = n9458_o[63:0];
  /* execute1.vhdl:468:35  */
  assign n9460_o = n9458_o[32];
  /* execute1.vhdl:468:49  */
  assign n9461_o = n9423_o[32];
  /* execute1.vhdl:468:40  */
  assign n9462_o = n9460_o ^ n9461_o;
  /* execute1.vhdl:468:62  */
  assign n9463_o = b_in[32];
  /* execute1.vhdl:468:54  */
  assign n9464_o = n9462_o ^ n9463_o;
  /* execute1.vhdl:469:35  */
  assign n9465_o = n9458_o[64];
  /* execute1.vhdl:470:37  */
  assign n9467_o = n9423_o[31];
  /* execute1.vhdl:470:47  */
  assign n9468_o = b_in[31];
  /* execute1.vhdl:470:77  */
  assign n9469_o = n9458_o[31];
  /* execute1.vhdl:197:20  */
  assign n9474_o = carry_32 ^ n9469_o;
  /* execute1.vhdl:197:46  */
  assign n9475_o = n9467_o ^ n9468_o;
  /* execute1.vhdl:197:35  */
  assign n9476_o = ~n9475_o;
  /* execute1.vhdl:197:31  */
  assign n9477_o = n9474_o & n9476_o;
  /* execute1.vhdl:471:37  */
  assign n9479_o = n9423_o[63];
  /* execute1.vhdl:471:47  */
  assign n9480_o = b_in[63];
  /* execute1.vhdl:471:77  */
  assign n9481_o = n9458_o[63];
  /* execute1.vhdl:197:20  */
  assign n9486_o = carry_64 ^ n9481_o;
  /* execute1.vhdl:197:46  */
  assign n9487_o = n9479_o ^ n9480_o;
  /* execute1.vhdl:197:35  */
  assign n9488_o = ~n9487_o;
  /* execute1.vhdl:197:31  */
  assign n9489_o = n9486_o & n9488_o;
  /* execute1.vhdl:476:17  */
  assign n9490_o = n9139_o[342];
  /* execute1.vhdl:477:21  */
  assign n9491_o = n9139_o[341];
  /* execute1.vhdl:478:30  */
  assign n9492_o = a_in[31];
  /* execute1.vhdl:479:30  */
  assign n9493_o = b_in[31];
  /* execute1.vhdl:481:30  */
  assign n9494_o = a_in[63];
  /* execute1.vhdl:482:30  */
  assign n9495_o = b_in[63];
  /* execute1.vhdl:477:13  */
  assign n9496_o = n9491_o ? n9492_o : n9494_o;
  /* execute1.vhdl:477:13  */
  assign n9497_o = n9491_o ? n9493_o : n9495_o;
  /* execute1.vhdl:476:9  */
  assign n9499_o = n9490_o ? n9496_o : 1'b0;
  /* execute1.vhdl:476:9  */
  assign n9502_o = n9490_o ? n9497_o : 1'b0;
  /* execute1.vhdl:486:18  */
  assign n9504_o = ~n9499_o;
  /* execute1.vhdl:489:21  */
  assign n9505_o = -a_in;
  /* execute1.vhdl:486:9  */
  assign n9506_o = n9504_o ? a_in : n9505_o;
  /* execute1.vhdl:491:18  */
  assign n9507_o = ~n9502_o;
  /* execute1.vhdl:494:21  */
  assign n9508_o = -b_in;
  /* execute1.vhdl:491:9  */
  assign n9509_o = n9507_o ? b_in : n9508_o;
  /* execute1.vhdl:498:40  */
  assign n9510_o = n9139_o[342];
  /* execute1.vhdl:499:39  */
  assign n9511_o = n9139_o[341];
  /* execute1.vhdl:502:17  */
  assign n9514_o = n9139_o[9:4];
  /* execute1.vhdl:502:27  */
  assign n9516_o = n9514_o == 6'b100101;
  /* execute1.vhdl:502:9  */
  assign n9518_o = n9516_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:507:21  */
  assign n9519_o = n9139_o[369];
  /* execute1.vhdl:507:26  */
  assign n9520_o = ~n9519_o;
  /* execute1.vhdl:510:21  */
  assign n9521_o = n9139_o[342];
  /* execute1.vhdl:511:57  */
  assign n9522_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9523_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9524_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9525_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9526_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9527_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9528_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9529_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9530_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9531_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9532_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9533_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9534_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9535_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9536_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9537_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9538_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9539_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9540_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9541_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9542_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9543_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9544_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9545_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9546_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9547_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9548_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9549_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9550_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9551_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9552_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9553_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9554_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9555_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9556_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9557_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9558_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9559_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9560_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9561_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9562_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9563_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9564_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9565_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9566_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9567_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9568_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9569_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9570_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9571_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9572_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9573_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9574_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9575_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9576_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9577_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9578_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9579_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9580_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9581_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9582_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9583_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9584_o = c_in[63];
  /* execute1.vhdl:511:57  */
  assign n9585_o = c_in[63];
  assign n9586_o = {n9522_o, n9523_o, n9524_o, n9525_o};
  assign n9587_o = {n9526_o, n9527_o, n9528_o, n9529_o};
  assign n9588_o = {n9530_o, n9531_o, n9532_o, n9533_o};
  assign n9589_o = {n9534_o, n9535_o, n9536_o, n9537_o};
  assign n9590_o = {n9538_o, n9539_o, n9540_o, n9541_o};
  assign n9591_o = {n9542_o, n9543_o, n9544_o, n9545_o};
  assign n9592_o = {n9546_o, n9547_o, n9548_o, n9549_o};
  assign n9593_o = {n9550_o, n9551_o, n9552_o, n9553_o};
  assign n9594_o = {n9554_o, n9555_o, n9556_o, n9557_o};
  assign n9595_o = {n9558_o, n9559_o, n9560_o, n9561_o};
  assign n9596_o = {n9562_o, n9563_o, n9564_o, n9565_o};
  assign n9597_o = {n9566_o, n9567_o, n9568_o, n9569_o};
  assign n9598_o = {n9570_o, n9571_o, n9572_o, n9573_o};
  assign n9599_o = {n9574_o, n9575_o, n9576_o, n9577_o};
  assign n9600_o = {n9578_o, n9579_o, n9580_o, n9581_o};
  assign n9601_o = {n9582_o, n9583_o, n9584_o, n9585_o};
  assign n9602_o = {n9586_o, n9587_o, n9588_o, n9589_o};
  assign n9603_o = {n9590_o, n9591_o, n9592_o, n9593_o};
  assign n9604_o = {n9594_o, n9595_o, n9596_o, n9597_o};
  assign n9605_o = {n9598_o, n9599_o, n9600_o, n9601_o};
  assign n9606_o = {n9602_o, n9603_o, n9604_o, n9605_o};
  /* execute1.vhdl:510:13  */
  assign n9608_o = n9521_o ? n9606_o : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  assign n9609_o = {n9608_o, c_in};
  /* execute1.vhdl:507:9  */
  assign n9611_o = n9520_o ? n9609_o : 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* execute1.vhdl:514:19  */
  assign n9613_o = n9499_o ^ n9502_o;
  /* execute1.vhdl:515:23  */
  assign n9614_o = ~n9611_o;
  /* execute1.vhdl:514:9  */
  assign n9615_o = n9613_o ? n9614_o : n9611_o;
  /* execute1.vhdl:518:40  */
  assign n9616_o = n9139_o[341];
  /* execute1.vhdl:519:43  */
  assign n9617_o = n9499_o ^ n9502_o;
  /* execute1.vhdl:521:74  */
  assign n9618_o = x_to_divider[132];
  /* execute1.vhdl:521:57  */
  assign n9619_o = ~n9618_o;
  /* execute1.vhdl:521:53  */
  assign n9620_o = n9502_o & n9619_o;
  /* execute1.vhdl:521:42  */
  assign n9621_o = n9499_o ^ n9620_o;
  /* execute1.vhdl:522:17  */
  assign n9622_o = n9139_o[341];
  /* execute1.vhdl:522:26  */
  assign n9623_o = ~n9622_o;
  /* execute1.vhdl:526:21  */
  assign n9624_o = n9139_o[9:4];
  /* execute1.vhdl:526:31  */
  assign n9626_o = n9624_o == 6'b010110;
  /* execute1.vhdl:526:13  */
  assign n9628_o = n9626_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:533:72  */
  assign n9629_o = n9506_o[31:0];
  /* execute1.vhdl:533:48  */
  assign n9631_o = {32'b00000000000000000000000000000000, n9629_o};
  /* execute1.vhdl:534:72  */
  assign n9632_o = n9509_o[31:0];
  /* execute1.vhdl:534:48  */
  assign n9634_o = {32'b00000000000000000000000000000000, n9632_o};
  /* execute1.vhdl:536:21  */
  assign n9636_o = n9139_o[9:4];
  /* execute1.vhdl:536:31  */
  assign n9638_o = n9636_o == 6'b010110;
  /* execute1.vhdl:537:64  */
  assign n9639_o = n9506_o[31:0];
  /* execute1.vhdl:537:79  */
  assign n9641_o = {n9639_o, 32'b00000000000000000000000000000000};
  /* execute1.vhdl:539:78  */
  assign n9642_o = n9506_o[31:0];
  /* execute1.vhdl:539:54  */
  assign n9644_o = {32'b00000000000000000000000000000000, n9642_o};
  /* execute1.vhdl:536:13  */
  assign n9645_o = n9638_o ? n9641_o : n9644_o;
  /* execute1.vhdl:541:73  */
  assign n9646_o = n9509_o[31:0];
  /* execute1.vhdl:541:49  */
  assign n9648_o = {32'b00000000000000000000000000000000, n9646_o};
  assign n9649_o = {n9634_o, n9631_o};
  assign n9650_o = {n9509_o, n9506_o};
  /* execute1.vhdl:522:9  */
  assign n9651_o = n9623_o ? n9650_o : n9649_o;
  assign n9652_o = {n9648_o, n9645_o};
  assign n9653_o = {n9509_o, n9506_o};
  /* execute1.vhdl:522:9  */
  assign n9654_o = n9623_o ? n9653_o : n9652_o;
  /* execute1.vhdl:522:9  */
  assign n9655_o = n9623_o ? n9628_o : 1'b0;
  /* execute1.vhdl:544:32  */
  assign n9656_o = current[388:387];
  /* execute1.vhdl:549:58  */
  assign n9657_o = multiply_to_x[64:1];
  /* execute1.vhdl:545:13  */
  assign n9659_o = n9656_o == 2'b00;
  /* execute1.vhdl:552:54  */
  assign n9660_o = multiply_to_x[128:65];
  /* execute1.vhdl:551:13  */
  assign n9662_o = n9656_o == 2'b01;
  /* execute1.vhdl:554:54  */
  assign n9663_o = multiply_to_x[64:33];
  /* execute1.vhdl:555:54  */
  assign n9664_o = multiply_to_x[64:33];
  /* execute1.vhdl:554:69  */
  assign n9665_o = {n9663_o, n9664_o};
  /* execute1.vhdl:553:13  */
  assign n9667_o = n9656_o == 2'b10;
  /* execute1.vhdl:557:47  */
  assign n9668_o = divider_to_x[64:1];
  assign n9669_o = {n9667_o, n9662_o, n9659_o};
  /* execute1.vhdl:544:9  */
  always @*
    case (n9669_o)
      3'b100: n9670_o = n9665_o;
      3'b010: n9670_o = n9660_o;
      3'b001: n9670_o = n9657_o;
      default: n9670_o = n9668_o;
    endcase
  /* execute1.vhdl:561:22  */
  assign n9671_o = current[389:387];
  /* execute1.vhdl:562:13  */
  assign n9673_o = n9671_o == 3'b000;
  /* execute1.vhdl:570:29  */
  assign n9674_o = a_in[4];
  /* execute1.vhdl:570:42  */
  assign n9675_o = b_in[4];
  /* execute1.vhdl:570:34  */
  assign n9676_o = n9674_o ^ n9675_o;
  /* execute1.vhdl:570:65  */
  assign n9677_o = n9458_o[4];
  /* execute1.vhdl:570:47  */
  assign n9678_o = n9676_o ^ n9677_o;
  /* execute1.vhdl:570:71  */
  assign n9679_o = ~n9678_o;
  /* execute1.vhdl:570:21  */
  assign n9682_o = n9679_o ? 4'b0110 : 4'b0000;
  /* execute1.vhdl:570:29  */
  assign n9685_o = a_in[8];
  /* execute1.vhdl:570:42  */
  assign n9686_o = b_in[8];
  /* execute1.vhdl:570:34  */
  assign n9687_o = n9685_o ^ n9686_o;
  /* execute1.vhdl:570:65  */
  assign n9688_o = n9458_o[8];
  /* execute1.vhdl:570:47  */
  assign n9689_o = n9687_o ^ n9688_o;
  /* execute1.vhdl:570:71  */
  assign n9690_o = ~n9689_o;
  assign n9692_o = n9683_o[7:4];
  /* execute1.vhdl:570:21  */
  assign n9693_o = n9690_o ? 4'b0110 : n9692_o;
  /* execute1.vhdl:570:29  */
  assign n9695_o = a_in[12];
  /* execute1.vhdl:570:42  */
  assign n9696_o = b_in[12];
  /* execute1.vhdl:570:34  */
  assign n9697_o = n9695_o ^ n9696_o;
  /* execute1.vhdl:570:65  */
  assign n9698_o = n9458_o[12];
  /* execute1.vhdl:570:47  */
  assign n9699_o = n9697_o ^ n9698_o;
  /* execute1.vhdl:570:71  */
  assign n9700_o = ~n9699_o;
  assign n9702_o = n9683_o[11:8];
  /* execute1.vhdl:570:21  */
  assign n9703_o = n9700_o ? 4'b0110 : n9702_o;
  /* execute1.vhdl:570:29  */
  assign n9705_o = a_in[16];
  /* execute1.vhdl:570:42  */
  assign n9706_o = b_in[16];
  /* execute1.vhdl:570:34  */
  assign n9707_o = n9705_o ^ n9706_o;
  /* execute1.vhdl:570:65  */
  assign n9708_o = n9458_o[16];
  /* execute1.vhdl:570:47  */
  assign n9709_o = n9707_o ^ n9708_o;
  /* execute1.vhdl:570:71  */
  assign n9710_o = ~n9709_o;
  assign n9712_o = n9683_o[15:12];
  /* execute1.vhdl:570:21  */
  assign n9713_o = n9710_o ? 4'b0110 : n9712_o;
  /* execute1.vhdl:570:29  */
  assign n9715_o = a_in[20];
  /* execute1.vhdl:570:42  */
  assign n9716_o = b_in[20];
  /* execute1.vhdl:570:34  */
  assign n9717_o = n9715_o ^ n9716_o;
  /* execute1.vhdl:570:65  */
  assign n9718_o = n9458_o[20];
  /* execute1.vhdl:570:47  */
  assign n9719_o = n9717_o ^ n9718_o;
  /* execute1.vhdl:570:71  */
  assign n9720_o = ~n9719_o;
  assign n9722_o = n9683_o[19:16];
  /* execute1.vhdl:570:21  */
  assign n9723_o = n9720_o ? 4'b0110 : n9722_o;
  /* execute1.vhdl:570:29  */
  assign n9725_o = a_in[24];
  /* execute1.vhdl:570:42  */
  assign n9726_o = b_in[24];
  /* execute1.vhdl:570:34  */
  assign n9727_o = n9725_o ^ n9726_o;
  /* execute1.vhdl:570:65  */
  assign n9728_o = n9458_o[24];
  /* execute1.vhdl:570:47  */
  assign n9729_o = n9727_o ^ n9728_o;
  /* execute1.vhdl:570:71  */
  assign n9730_o = ~n9729_o;
  assign n9732_o = n9683_o[23:20];
  /* execute1.vhdl:570:21  */
  assign n9733_o = n9730_o ? 4'b0110 : n9732_o;
  /* execute1.vhdl:570:29  */
  assign n9735_o = a_in[28];
  /* execute1.vhdl:570:42  */
  assign n9736_o = b_in[28];
  /* execute1.vhdl:570:34  */
  assign n9737_o = n9735_o ^ n9736_o;
  /* execute1.vhdl:570:65  */
  assign n9738_o = n9458_o[28];
  /* execute1.vhdl:570:47  */
  assign n9739_o = n9737_o ^ n9738_o;
  /* execute1.vhdl:570:71  */
  assign n9740_o = ~n9739_o;
  assign n9742_o = n9683_o[27:24];
  /* execute1.vhdl:570:21  */
  assign n9743_o = n9740_o ? 4'b0110 : n9742_o;
  /* execute1.vhdl:570:29  */
  assign n9745_o = a_in[32];
  /* execute1.vhdl:570:42  */
  assign n9746_o = b_in[32];
  /* execute1.vhdl:570:34  */
  assign n9747_o = n9745_o ^ n9746_o;
  /* execute1.vhdl:570:65  */
  assign n9748_o = n9458_o[32];
  /* execute1.vhdl:570:47  */
  assign n9749_o = n9747_o ^ n9748_o;
  /* execute1.vhdl:570:71  */
  assign n9750_o = ~n9749_o;
  assign n9752_o = n9683_o[31:28];
  /* execute1.vhdl:570:21  */
  assign n9753_o = n9750_o ? 4'b0110 : n9752_o;
  /* execute1.vhdl:570:29  */
  assign n9755_o = a_in[36];
  /* execute1.vhdl:570:42  */
  assign n9756_o = b_in[36];
  /* execute1.vhdl:570:34  */
  assign n9757_o = n9755_o ^ n9756_o;
  /* execute1.vhdl:570:65  */
  assign n9758_o = n9458_o[36];
  /* execute1.vhdl:570:47  */
  assign n9759_o = n9757_o ^ n9758_o;
  /* execute1.vhdl:570:71  */
  assign n9760_o = ~n9759_o;
  assign n9762_o = n9683_o[35:32];
  /* execute1.vhdl:570:21  */
  assign n9763_o = n9760_o ? 4'b0110 : n9762_o;
  /* execute1.vhdl:570:29  */
  assign n9765_o = a_in[40];
  /* execute1.vhdl:570:42  */
  assign n9766_o = b_in[40];
  /* execute1.vhdl:570:34  */
  assign n9767_o = n9765_o ^ n9766_o;
  /* execute1.vhdl:570:65  */
  assign n9768_o = n9458_o[40];
  /* execute1.vhdl:570:47  */
  assign n9769_o = n9767_o ^ n9768_o;
  /* execute1.vhdl:570:71  */
  assign n9770_o = ~n9769_o;
  assign n9772_o = n9683_o[39:36];
  /* execute1.vhdl:570:21  */
  assign n9773_o = n9770_o ? 4'b0110 : n9772_o;
  /* execute1.vhdl:570:29  */
  assign n9775_o = a_in[44];
  /* execute1.vhdl:570:42  */
  assign n9776_o = b_in[44];
  /* execute1.vhdl:570:34  */
  assign n9777_o = n9775_o ^ n9776_o;
  /* execute1.vhdl:570:65  */
  assign n9778_o = n9458_o[44];
  /* execute1.vhdl:570:47  */
  assign n9779_o = n9777_o ^ n9778_o;
  /* execute1.vhdl:570:71  */
  assign n9780_o = ~n9779_o;
  assign n9782_o = n9683_o[43:40];
  /* execute1.vhdl:570:21  */
  assign n9783_o = n9780_o ? 4'b0110 : n9782_o;
  /* execute1.vhdl:570:29  */
  assign n9785_o = a_in[48];
  /* execute1.vhdl:570:42  */
  assign n9786_o = b_in[48];
  /* execute1.vhdl:570:34  */
  assign n9787_o = n9785_o ^ n9786_o;
  /* execute1.vhdl:570:65  */
  assign n9788_o = n9458_o[48];
  /* execute1.vhdl:570:47  */
  assign n9789_o = n9787_o ^ n9788_o;
  /* execute1.vhdl:570:71  */
  assign n9790_o = ~n9789_o;
  assign n9792_o = n9683_o[47:44];
  /* execute1.vhdl:570:21  */
  assign n9793_o = n9790_o ? 4'b0110 : n9792_o;
  /* execute1.vhdl:570:29  */
  assign n9795_o = a_in[52];
  /* execute1.vhdl:570:42  */
  assign n9796_o = b_in[52];
  /* execute1.vhdl:570:34  */
  assign n9797_o = n9795_o ^ n9796_o;
  /* execute1.vhdl:570:65  */
  assign n9798_o = n9458_o[52];
  /* execute1.vhdl:570:47  */
  assign n9799_o = n9797_o ^ n9798_o;
  /* execute1.vhdl:570:71  */
  assign n9800_o = ~n9799_o;
  assign n9802_o = n9683_o[51:48];
  /* execute1.vhdl:570:21  */
  assign n9803_o = n9800_o ? 4'b0110 : n9802_o;
  /* execute1.vhdl:570:29  */
  assign n9805_o = a_in[56];
  /* execute1.vhdl:570:42  */
  assign n9806_o = b_in[56];
  /* execute1.vhdl:570:34  */
  assign n9807_o = n9805_o ^ n9806_o;
  /* execute1.vhdl:570:65  */
  assign n9808_o = n9458_o[56];
  /* execute1.vhdl:570:47  */
  assign n9809_o = n9807_o ^ n9808_o;
  /* execute1.vhdl:570:71  */
  assign n9810_o = ~n9809_o;
  assign n9812_o = n9683_o[55:52];
  /* execute1.vhdl:570:21  */
  assign n9813_o = n9810_o ? 4'b0110 : n9812_o;
  /* execute1.vhdl:570:29  */
  assign n9815_o = a_in[60];
  /* execute1.vhdl:570:42  */
  assign n9816_o = b_in[60];
  /* execute1.vhdl:570:34  */
  assign n9817_o = n9815_o ^ n9816_o;
  /* execute1.vhdl:570:65  */
  assign n9818_o = n9458_o[60];
  /* execute1.vhdl:570:47  */
  assign n9819_o = n9817_o ^ n9818_o;
  /* execute1.vhdl:570:71  */
  assign n9820_o = ~n9819_o;
  assign n9822_o = n9683_o[59:56];
  /* execute1.vhdl:570:21  */
  assign n9823_o = n9820_o ? 4'b0110 : n9822_o;
  assign n9824_o = n9683_o[63:60];
  /* execute1.vhdl:574:34  */
  assign n9825_o = n9458_o[64];
  /* execute1.vhdl:574:39  */
  assign n9826_o = ~n9825_o;
  /* execute1.vhdl:574:17  */
  assign n9828_o = n9826_o ? 4'b0110 : n9824_o;
  assign n9829_o = {n9828_o, n9823_o, n9813_o, n9803_o, n9793_o, n9783_o, n9773_o, n9763_o, n9753_o, n9743_o, n9733_o, n9723_o, n9713_o, n9703_o, n9693_o, n9682_o};
  /* execute1.vhdl:564:13  */
  assign n9831_o = n9671_o == 3'b001;
  /* execute1.vhdl:580:59  */
  assign n9833_o = n9139_o[374:343];
  /* insn_helpers.vhdl:211:23  */
  assign n9838_o = n9833_o[10:6];
  /* execute1.vhdl:581:28  */
  assign n9840_o = {27'b0, n9838_o};  //  uext
  /* execute1.vhdl:581:28  */
  assign n9842_o = 32'b00000000000000000000000000011111 - n9840_o;
  /* execute1.vhdl:581:28  */
  assign n9843_o = n9842_o[4:0];  // trunc
  /* execute1.vhdl:581:17  */
  assign n9846_o = n12615_o ? a_in : b_in;
  /* execute1.vhdl:578:13  */
  assign n9848_o = n9671_o == 3'b010;
  /* execute1.vhdl:590:31  */
  assign n9849_o = ~random_err;
  /* execute1.vhdl:591:35  */
  assign n9850_o = n9139_o[360:359];
  /* execute1.vhdl:593:62  */
  assign n9851_o = random_cond[31:0];
  /* execute1.vhdl:593:49  */
  assign n9853_o = {32'b00000000000000000000000000000000, n9851_o};
  /* execute1.vhdl:592:25  */
  assign n9855_o = n9850_o == 2'b00;
  /* execute1.vhdl:594:25  */
  assign n9857_o = n9850_o == 2'b10;
  assign n9858_o = {n9857_o, n9855_o};
  /* execute1.vhdl:591:21  */
  always @*
    case (n9858_o)
      2'b10: n9859_o = random_raw;
      2'b01: n9859_o = n9853_o;
      default: n9859_o = random_cond;
    endcase
  /* execute1.vhdl:590:17  */
  assign n9861_o = n9849_o ? n9859_o : 64'b1111111111111111111111111111111111111111111111111111111111111111;
  /* execute1.vhdl:587:13  */
  assign n9864_o = n9671_o == 3'b011;
  /* execute1.vhdl:603:37  */
  assign n9865_o = ctrl[191:128];
  /* execute1.vhdl:601:13  */
  assign n9867_o = n9671_o == 3'b100;
  /* execute1.vhdl:605:29  */
  assign n9868_o = n9139_o[363];
  /* execute1.vhdl:605:34  */
  assign n9869_o = ~n9868_o;
  /* execute1.vhdl:607:48  */
  assign n9871_o = {32'b00000000000000000000000000000000, cr_in};
  /* execute1.vhdl:610:55  */
  assign n9874_o = n9139_o[374:343];
  /* insn_helpers.vhdl:166:23  */
  assign n9879_o = n9874_o[19:12];
  /* crhelpers.vhdl:23:19  */
  assign n9884_o = n9879_o[7];
  /* crhelpers.vhdl:23:13  */
  assign n9888_o = n9884_o ? 1'b0 : 1'b1;
  /* crhelpers.vhdl:23:13  */
  assign n9892_o = n9884_o ? 1'b0 : 1'b1;
  /* crhelpers.vhdl:23:13  */
  assign n9894_o = n9884_o ? 3'b000 : 3'bX;
  /* crhelpers.vhdl:23:19  */
  assign n9895_o = n9879_o[6];
  /* crhelpers.vhdl:23:13  */
  assign n9898_o = n9905_o ? 1'b0 : n9888_o;
  /* crhelpers.vhdl:23:13  */
  assign n9900_o = n9906_o ? 1'b0 : n9892_o;
  /* crhelpers.vhdl:23:13  */
  assign n9901_o = n9907_o ? 3'b001 : n9894_o;
  /* crhelpers.vhdl:23:13  */
  assign n9902_o = n9895_o & n9888_o;
  /* crhelpers.vhdl:23:13  */
  assign n9903_o = n9895_o & n9888_o;
  /* crhelpers.vhdl:23:13  */
  assign n9904_o = n9895_o & n9888_o;
  /* crhelpers.vhdl:23:13  */
  assign n9905_o = n9888_o & n9902_o;
  /* crhelpers.vhdl:23:13  */
  assign n9906_o = n9888_o & n9903_o;
  /* crhelpers.vhdl:23:13  */
  assign n9907_o = n9888_o & n9904_o;
  /* crhelpers.vhdl:23:19  */
  assign n9908_o = n9879_o[5];
  /* crhelpers.vhdl:23:13  */
  assign n9911_o = n9918_o ? 1'b0 : n9898_o;
  /* crhelpers.vhdl:23:13  */
  assign n9913_o = n9919_o ? 1'b0 : n9900_o;
  /* crhelpers.vhdl:23:13  */
  assign n9914_o = n9920_o ? 3'b010 : n9901_o;
  /* crhelpers.vhdl:23:13  */
  assign n9915_o = n9908_o & n9898_o;
  /* crhelpers.vhdl:23:13  */
  assign n9916_o = n9908_o & n9898_o;
  /* crhelpers.vhdl:23:13  */
  assign n9917_o = n9908_o & n9898_o;
  /* crhelpers.vhdl:23:13  */
  assign n9918_o = n9898_o & n9915_o;
  /* crhelpers.vhdl:23:13  */
  assign n9919_o = n9898_o & n9916_o;
  /* crhelpers.vhdl:23:13  */
  assign n9920_o = n9898_o & n9917_o;
  /* crhelpers.vhdl:23:19  */
  assign n9921_o = n9879_o[4];
  /* crhelpers.vhdl:23:13  */
  assign n9924_o = n9931_o ? 1'b0 : n9911_o;
  /* crhelpers.vhdl:23:13  */
  assign n9926_o = n9932_o ? 1'b0 : n9913_o;
  /* crhelpers.vhdl:23:13  */
  assign n9927_o = n9933_o ? 3'b011 : n9914_o;
  /* crhelpers.vhdl:23:13  */
  assign n9928_o = n9921_o & n9911_o;
  /* crhelpers.vhdl:23:13  */
  assign n9929_o = n9921_o & n9911_o;
  /* crhelpers.vhdl:23:13  */
  assign n9930_o = n9921_o & n9911_o;
  /* crhelpers.vhdl:23:13  */
  assign n9931_o = n9911_o & n9928_o;
  /* crhelpers.vhdl:23:13  */
  assign n9932_o = n9911_o & n9929_o;
  /* crhelpers.vhdl:23:13  */
  assign n9933_o = n9911_o & n9930_o;
  /* crhelpers.vhdl:23:19  */
  assign n9934_o = n9879_o[3];
  /* crhelpers.vhdl:23:13  */
  assign n9937_o = n9944_o ? 1'b0 : n9924_o;
  /* crhelpers.vhdl:23:13  */
  assign n9939_o = n9945_o ? 1'b0 : n9926_o;
  /* crhelpers.vhdl:23:13  */
  assign n9940_o = n9946_o ? 3'b100 : n9927_o;
  /* crhelpers.vhdl:23:13  */
  assign n9941_o = n9934_o & n9924_o;
  /* crhelpers.vhdl:23:13  */
  assign n9942_o = n9934_o & n9924_o;
  /* crhelpers.vhdl:23:13  */
  assign n9943_o = n9934_o & n9924_o;
  /* crhelpers.vhdl:23:13  */
  assign n9944_o = n9924_o & n9941_o;
  /* crhelpers.vhdl:23:13  */
  assign n9945_o = n9924_o & n9942_o;
  /* crhelpers.vhdl:23:13  */
  assign n9946_o = n9924_o & n9943_o;
  /* crhelpers.vhdl:23:19  */
  assign n9947_o = n9879_o[2];
  /* crhelpers.vhdl:23:13  */
  assign n9950_o = n9957_o ? 1'b0 : n9937_o;
  /* crhelpers.vhdl:23:13  */
  assign n9952_o = n9958_o ? 1'b0 : n9939_o;
  /* crhelpers.vhdl:23:13  */
  assign n9953_o = n9959_o ? 3'b101 : n9940_o;
  /* crhelpers.vhdl:23:13  */
  assign n9954_o = n9947_o & n9937_o;
  /* crhelpers.vhdl:23:13  */
  assign n9955_o = n9947_o & n9937_o;
  /* crhelpers.vhdl:23:13  */
  assign n9956_o = n9947_o & n9937_o;
  /* crhelpers.vhdl:23:13  */
  assign n9957_o = n9937_o & n9954_o;
  /* crhelpers.vhdl:23:13  */
  assign n9958_o = n9937_o & n9955_o;
  /* crhelpers.vhdl:23:13  */
  assign n9959_o = n9937_o & n9956_o;
  /* crhelpers.vhdl:23:19  */
  assign n9960_o = n9879_o[1];
  /* crhelpers.vhdl:23:13  */
  assign n9963_o = n9970_o ? 1'b0 : n9950_o;
  /* crhelpers.vhdl:23:13  */
  assign n9965_o = n9971_o ? 1'b0 : n9952_o;
  /* crhelpers.vhdl:23:13  */
  assign n9966_o = n9972_o ? 3'b110 : n9953_o;
  /* crhelpers.vhdl:23:13  */
  assign n9967_o = n9960_o & n9950_o;
  /* crhelpers.vhdl:23:13  */
  assign n9968_o = n9960_o & n9950_o;
  /* crhelpers.vhdl:23:13  */
  assign n9969_o = n9960_o & n9950_o;
  /* crhelpers.vhdl:23:13  */
  assign n9970_o = n9950_o & n9967_o;
  /* crhelpers.vhdl:23:13  */
  assign n9971_o = n9950_o & n9968_o;
  /* crhelpers.vhdl:23:13  */
  assign n9972_o = n9950_o & n9969_o;
  /* crhelpers.vhdl:23:19  */
  assign n9973_o = n9879_o[0];
  /* crhelpers.vhdl:23:13  */
  assign n9978_o = n9984_o ? 1'b0 : n9965_o;
  /* crhelpers.vhdl:23:13  */
  assign n9979_o = n9985_o ? 3'b111 : n9966_o;
  /* crhelpers.vhdl:23:13  */
  assign n9981_o = n9973_o & n9963_o;
  /* crhelpers.vhdl:23:13  */
  assign n9982_o = n9973_o & n9963_o;
  /* crhelpers.vhdl:23:13  */
  assign n9984_o = n9963_o & n9981_o;
  /* crhelpers.vhdl:23:13  */
  assign n9985_o = n9963_o & n9982_o;
  /* crhelpers.vhdl:30:9  */
  assign n9991_o = n9978_o ? 3'b111 : n9979_o;
  /* execute1.vhdl:615:34  */
  assign n9992_o = {29'b0, n9991_o};  //  uext
  /* execute1.vhdl:615:34  */
  assign n9994_o = n9992_o == 32'b00000000000000000000000000000000;
  /* execute1.vhdl:616:63  */
  assign n9995_o = cr_in[31:28];
  /* execute1.vhdl:615:25  */
  assign n9997_o = n9994_o ? n9995_o : 4'b0000;
  assign n9999_o = n9998_o[63:32];
  /* execute1.vhdl:615:34  */
  assign n10001_o = {29'b0, n9991_o};  //  uext
  /* execute1.vhdl:615:34  */
  assign n10003_o = n10001_o == 32'b00000000000000000000000000000001;
  /* execute1.vhdl:616:63  */
  assign n10004_o = cr_in[27:24];
  assign n10005_o = n9998_o[27:24];
  /* execute1.vhdl:615:25  */
  assign n10006_o = n10003_o ? n10004_o : n10005_o;
  /* execute1.vhdl:615:34  */
  assign n10008_o = {29'b0, n9991_o};  //  uext
  /* execute1.vhdl:615:34  */
  assign n10010_o = n10008_o == 32'b00000000000000000000000000000010;
  /* execute1.vhdl:616:63  */
  assign n10011_o = cr_in[23:20];
  assign n10012_o = n9998_o[23:20];
  /* execute1.vhdl:615:25  */
  assign n10013_o = n10010_o ? n10011_o : n10012_o;
  /* execute1.vhdl:615:34  */
  assign n10015_o = {29'b0, n9991_o};  //  uext
  /* execute1.vhdl:615:34  */
  assign n10017_o = n10015_o == 32'b00000000000000000000000000000011;
  /* execute1.vhdl:616:63  */
  assign n10018_o = cr_in[19:16];
  assign n10019_o = n9998_o[19:16];
  /* execute1.vhdl:615:25  */
  assign n10020_o = n10017_o ? n10018_o : n10019_o;
  /* execute1.vhdl:615:34  */
  assign n10022_o = {29'b0, n9991_o};  //  uext
  /* execute1.vhdl:615:34  */
  assign n10024_o = n10022_o == 32'b00000000000000000000000000000100;
  /* execute1.vhdl:616:63  */
  assign n10025_o = cr_in[15:12];
  assign n10026_o = n9998_o[15:12];
  /* execute1.vhdl:615:25  */
  assign n10027_o = n10024_o ? n10025_o : n10026_o;
  /* execute1.vhdl:615:34  */
  assign n10029_o = {29'b0, n9991_o};  //  uext
  /* execute1.vhdl:615:34  */
  assign n10031_o = n10029_o == 32'b00000000000000000000000000000101;
  /* execute1.vhdl:616:63  */
  assign n10032_o = cr_in[11:8];
  assign n10033_o = n9998_o[11:8];
  /* execute1.vhdl:615:25  */
  assign n10034_o = n10031_o ? n10032_o : n10033_o;
  /* execute1.vhdl:615:34  */
  assign n10036_o = {29'b0, n9991_o};  //  uext
  /* execute1.vhdl:615:34  */
  assign n10038_o = n10036_o == 32'b00000000000000000000000000000110;
  /* execute1.vhdl:616:63  */
  assign n10039_o = cr_in[7:4];
  assign n10040_o = n9998_o[7:4];
  /* execute1.vhdl:615:25  */
  assign n10041_o = n10038_o ? n10039_o : n10040_o;
  assign n10042_o = n9998_o[3:0];
  /* execute1.vhdl:615:34  */
  assign n10043_o = {29'b0, n9991_o};  //  uext
  /* execute1.vhdl:615:34  */
  assign n10045_o = n10043_o == 32'b00000000000000000000000000000111;
  /* execute1.vhdl:616:63  */
  assign n10046_o = cr_in[3:0];
  /* execute1.vhdl:615:25  */
  assign n10047_o = n10045_o ? n10046_o : n10042_o;
  assign n10048_o = {n9999_o, n9997_o, n10006_o, n10013_o, n10020_o, n10027_o, n10034_o, n10041_o, n10047_o};
  /* execute1.vhdl:605:17  */
  assign n10049_o = n9869_o ? n9871_o : n10048_o;
  /* execute1.vhdl:604:13  */
  assign n10056_o = n9671_o == 3'b101;
  /* execute1.vhdl:623:38  */
  assign n10058_o = n9139_o[374:343];
  /* insn_helpers.vhdl:141:23  */
  assign n10063_o = n10058_o[20:18];
  /* execute1.vhdl:624:26  */
  assign n10064_o = {28'b0, n10063_o};  //  uext
  /* execute1.vhdl:624:52  */
  assign n10065_o = {1'b0, n10064_o};  //  uext
  /* execute1.vhdl:624:52  */
  assign n10067_o = n10065_o * 32'b00000000000000000000000000000100; // smul
  /* execute1.vhdl:624:17  */
  assign n10068_o = n10067_o[4:0];  // trunc
  /* execute1.vhdl:626:29  */
  assign n10069_o = {27'b0, n10068_o};  //  uext
  /* execute1.vhdl:626:29  */
  assign n10071_o = 32'b00000000000000000000000000011111 - n10069_o;
  /* execute1.vhdl:626:29  */
  assign n10072_o = n10071_o[4:0];  // trunc
  /* execute1.vhdl:628:32  */
  assign n10075_o = {27'b0, n10068_o};  //  uext
  /* execute1.vhdl:628:32  */
  assign n10077_o = 32'b00000000000000000000000000011110 - n10075_o;
  /* execute1.vhdl:628:32  */
  assign n10078_o = n10077_o[4:0];  // trunc
  /* execute1.vhdl:628:17  */
  assign n10083_o = n12723_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:626:17  */
  assign n10085_o = n12669_o ? 1'b1 : n10083_o;
  /* execute1.vhdl:626:17  */
  assign n10088_o = n12669_o ? 63'b111111111111111111111111111111111111111111111111111111111111111 : 63'b000000000000000000000000000000000000000000000000000000000000000;
  assign n10091_o = {n10088_o, n10085_o};
  /* execute1.vhdl:621:13  */
  assign n10093_o = n9671_o == 3'b110;
  assign n10094_o = {n10093_o, n10056_o, n9867_o, n9864_o, n9848_o, n9831_o, n9673_o};
  /* execute1.vhdl:561:9  */
  always @*
    case (n10094_o)
      7'b1000000: n10097_o = n10091_o;
      7'b0100000: n10097_o = n10049_o;
      7'b0010000: n10097_o = n9865_o;
      7'b0001000: n10097_o = n9861_o;
      7'b0000100: n10097_o = n9846_o;
      7'b0000010: n10097_o = n9829_o;
      7'b0000001: n10097_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      default: n10097_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* execute1.vhdl:638:17  */
  assign n10144_o = n9139_o[9:4];
  /* execute1.vhdl:638:27  */
  assign n10146_o = n10144_o == 6'b001001;
  /* execute1.vhdl:639:30  */
  assign n10148_o = n9139_o[374:343];
  /* insn_helpers.vhdl:86:23  */
  assign n10153_o = n10148_o[21];
  /* execute1.vhdl:641:27  */
  assign n10154_o = n9139_o[341];
  /* execute1.vhdl:641:18  */
  assign n10155_o = ~n10154_o;
  /* execute1.vhdl:638:9  */
  assign n10156_o = n10146_o ? n10153_o : n10155_o;
  /* execute1.vhdl:643:32  */
  assign n10157_o = a_in[31:0];
  /* execute1.vhdl:643:54  */
  assign n10158_o = b_in[31:0];
  /* execute1.vhdl:643:46  */
  assign n10159_o = n10157_o ^ n10158_o;
  /* execute1.vhdl:643:24  */
  assign n10160_o = |(n10159_o);
  /* execute1.vhdl:643:19  */
  assign n10161_o = ~n10160_o;
  /* execute1.vhdl:644:32  */
  assign n10162_o = a_in[63:32];
  /* execute1.vhdl:644:55  */
  assign n10163_o = b_in[63:32];
  /* execute1.vhdl:644:47  */
  assign n10164_o = n10162_o ^ n10163_o;
  /* execute1.vhdl:644:24  */
  assign n10165_o = |(n10164_o);
  /* execute1.vhdl:644:19  */
  assign n10166_o = ~n10165_o;
  /* execute1.vhdl:645:32  */
  assign n10167_o = ~n10156_o;
  /* execute1.vhdl:645:38  */
  assign n10168_o = n10167_o | n10166_o;
  /* execute1.vhdl:645:25  */
  assign n10169_o = n10161_o & n10168_o;
  /* execute1.vhdl:651:29  */
  assign n10170_o = a_in[30:0];
  /* execute1.vhdl:651:59  */
  assign n10171_o = b_in[30:0];
  /* execute1.vhdl:651:44  */
  assign n10172_o = $unsigned(n10170_o) < $unsigned(n10171_o);
  /* execute1.vhdl:651:13  */
  assign n10175_o = n10172_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:654:29  */
  assign n10177_o = a_in[62:31];
  /* execute1.vhdl:654:60  */
  assign n10178_o = b_in[62:31];
  /* execute1.vhdl:654:45  */
  assign n10179_o = $unsigned(n10177_o) < $unsigned(n10178_o);
  /* execute1.vhdl:654:13  */
  assign n10182_o = n10179_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:659:30  */
  assign n10184_o = a_in[63];
  /* execute1.vhdl:660:30  */
  assign n10185_o = b_in[63];
  /* execute1.vhdl:661:53  */
  assign n10186_o = a_in[31];
  /* execute1.vhdl:661:67  */
  assign n10187_o = b_in[31];
  /* execute1.vhdl:661:58  */
  assign n10188_o = ~(n10186_o ^ n10187_o);
  /* execute1.vhdl:661:44  */
  assign n10189_o = n10166_o & n10188_o;
  /* execute1.vhdl:661:73  */
  assign n10190_o = n10189_o & n10175_o;
  /* execute1.vhdl:661:33  */
  assign n10191_o = n10182_o | n10190_o;
  /* execute1.vhdl:664:30  */
  assign n10192_o = a_in[31];
  /* execute1.vhdl:665:30  */
  assign n10193_o = b_in[31];
  /* execute1.vhdl:657:13  */
  assign n10194_o = n10156_o ? n10184_o : n10192_o;
  /* execute1.vhdl:657:13  */
  assign n10195_o = n10156_o ? n10185_o : n10193_o;
  /* execute1.vhdl:657:13  */
  assign n10196_o = n10156_o ? n10191_o : n10175_o;
  /* execute1.vhdl:668:22  */
  assign n10197_o = n10194_o != n10195_o;
  /* execute1.vhdl:671:34  */
  assign n10198_o = {n10194_o, n10195_o};
  /* execute1.vhdl:671:42  */
  assign n10200_o = {n10198_o, 1'b0};
  /* execute1.vhdl:671:48  */
  assign n10201_o = {n10200_o, n10195_o};
  /* execute1.vhdl:671:56  */
  assign n10202_o = {n10201_o, n10194_o};
  /* execute1.vhdl:675:35  */
  assign n10203_o = ~n10196_o;
  /* execute1.vhdl:675:33  */
  assign n10204_o = {n10196_o, n10203_o};
  /* execute1.vhdl:675:44  */
  assign n10206_o = {n10204_o, 1'b0};
  /* execute1.vhdl:675:50  */
  assign n10207_o = {n10206_o, n10196_o};
  /* execute1.vhdl:675:59  */
  assign n10208_o = ~n10196_o;
  /* execute1.vhdl:675:57  */
  assign n10209_o = {n10207_o, n10208_o};
  /* execute1.vhdl:668:13  */
  assign n10210_o = n10197_o ? n10202_o : n10209_o;
  /* execute1.vhdl:645:9  */
  assign n10212_o = n10169_o ? 5'b00100 : n10210_o;
  /* execute1.vhdl:680:28  */
  assign n10219_o = n9139_o[374:343];
  /* insn_helpers.vhdl:136:23  */
  assign n10224_o = n10219_o[25:23];
  /* execute1.vhdl:683:22  */
  assign n10226_o = current[389:387];
  /* execute1.vhdl:686:25  */
  assign n10227_o = n9139_o[342];
  /* execute1.vhdl:687:38  */
  assign n10228_o = trapval[4:2];
  /* execute1.vhdl:687:61  */
  assign n10229_o = xerc_in[4];
  /* execute1.vhdl:687:51  */
  assign n10230_o = {n10228_o, n10229_o};
  /* execute1.vhdl:689:38  */
  assign n10231_o = trapval[1:0];
  /* execute1.vhdl:689:60  */
  assign n10232_o = trapval[2];
  /* execute1.vhdl:689:51  */
  assign n10233_o = {n10231_o, n10232_o};
  /* execute1.vhdl:689:74  */
  assign n10234_o = xerc_in[4];
  /* execute1.vhdl:689:64  */
  assign n10235_o = {n10233_o, n10234_o};
  /* execute1.vhdl:686:17  */
  assign n10236_o = n10227_o ? n10230_o : n10235_o;
  /* execute1.vhdl:684:13  */
  assign n10238_o = n10226_o == 3'b000;
  /* execute1.vhdl:692:61  */
  assign n10241_o = n9139_o[374:343];
  /* insn_helpers.vhdl:86:23  */
  assign n10246_o = n10241_o[21];
  /* ppc_fx_insns.vhdl:770:29  */
  assign n10253_o = a_in[7:0];
  /* ppc_fx_insns.vhdl:771:32  */
  assign n10255_o = b_in[7:0];
  /* ppc_fx_insns.vhdl:771:18  */
  assign n10256_o = $unsigned(n10253_o) >= $unsigned(n10255_o);
  /* ppc_fx_insns.vhdl:771:66  */
  assign n10257_o = b_in[15:8];
  /* ppc_fx_insns.vhdl:771:52  */
  assign n10258_o = $unsigned(n10253_o) <= $unsigned(n10257_o);
  /* ppc_fx_insns.vhdl:771:46  */
  assign n10259_o = n10256_o & n10258_o;
  /* ppc_fx_insns.vhdl:773:47  */
  assign n10260_o = b_in[23:16];
  /* ppc_fx_insns.vhdl:773:33  */
  assign n10261_o = $unsigned(n10253_o) >= $unsigned(n10260_o);
  /* ppc_fx_insns.vhdl:773:27  */
  assign n10262_o = n10246_o & n10261_o;
  /* ppc_fx_insns.vhdl:773:83  */
  assign n10263_o = b_in[31:24];
  /* ppc_fx_insns.vhdl:773:69  */
  assign n10264_o = $unsigned(n10253_o) <= $unsigned(n10263_o);
  /* ppc_fx_insns.vhdl:773:63  */
  assign n10265_o = n10262_o & n10264_o;
  /* ppc_fx_insns.vhdl:773:13  */
  assign n10268_o = n10265_o ? 1'b1 : 1'b0;
  /* ppc_fx_insns.vhdl:771:13  */
  assign n10270_o = n10259_o ? 1'b1 : n10268_o;
  /* ppc_fx_insns.vhdl:776:24  */
  assign n10273_o = {1'b0, n10270_o};
  /* ppc_fx_insns.vhdl:776:32  */
  assign n10275_o = {n10273_o, 2'b00};
  /* execute1.vhdl:691:13  */
  assign n10277_o = n10226_o == 3'b001;
  /* ppc_fx_insns.vhdl:758:22  */
  assign n10285_o = a_in[7:0];
  /* ppc_fx_insns.vhdl:758:39  */
  assign n10286_o = b_in[7:0];
  /* ppc_fx_insns.vhdl:758:35  */
  assign n10287_o = n10285_o == n10286_o;
  /* ppc_fx_insns.vhdl:758:17  */
  assign n10290_o = n10287_o ? 1'b1 : 1'b0;
  /* ppc_fx_insns.vhdl:758:22  */
  assign n10292_o = a_in[7:0];
  /* ppc_fx_insns.vhdl:758:39  */
  assign n10293_o = b_in[15:8];
  /* ppc_fx_insns.vhdl:758:35  */
  assign n10294_o = n10292_o == n10293_o;
  /* ppc_fx_insns.vhdl:758:17  */
  assign n10296_o = n10294_o ? 1'b1 : n10290_o;
  /* ppc_fx_insns.vhdl:758:22  */
  assign n10297_o = a_in[7:0];
  /* ppc_fx_insns.vhdl:758:39  */
  assign n10298_o = b_in[23:16];
  /* ppc_fx_insns.vhdl:758:35  */
  assign n10299_o = n10297_o == n10298_o;
  /* ppc_fx_insns.vhdl:758:17  */
  assign n10301_o = n10299_o ? 1'b1 : n10296_o;
  /* ppc_fx_insns.vhdl:758:22  */
  assign n10302_o = a_in[7:0];
  /* ppc_fx_insns.vhdl:758:39  */
  assign n10303_o = b_in[31:24];
  /* ppc_fx_insns.vhdl:758:35  */
  assign n10304_o = n10302_o == n10303_o;
  /* ppc_fx_insns.vhdl:758:17  */
  assign n10306_o = n10304_o ? 1'b1 : n10301_o;
  /* ppc_fx_insns.vhdl:758:22  */
  assign n10307_o = a_in[7:0];
  /* ppc_fx_insns.vhdl:758:39  */
  assign n10308_o = b_in[39:32];
  /* ppc_fx_insns.vhdl:758:35  */
  assign n10309_o = n10307_o == n10308_o;
  /* ppc_fx_insns.vhdl:758:17  */
  assign n10311_o = n10309_o ? 1'b1 : n10306_o;
  /* ppc_fx_insns.vhdl:758:22  */
  assign n10312_o = a_in[7:0];
  /* ppc_fx_insns.vhdl:758:39  */
  assign n10313_o = b_in[47:40];
  /* ppc_fx_insns.vhdl:758:35  */
  assign n10314_o = n10312_o == n10313_o;
  /* ppc_fx_insns.vhdl:758:17  */
  assign n10316_o = n10314_o ? 1'b1 : n10311_o;
  /* ppc_fx_insns.vhdl:758:22  */
  assign n10317_o = a_in[7:0];
  /* ppc_fx_insns.vhdl:758:39  */
  assign n10318_o = b_in[55:48];
  /* ppc_fx_insns.vhdl:758:35  */
  assign n10319_o = n10317_o == n10318_o;
  /* ppc_fx_insns.vhdl:758:17  */
  assign n10321_o = n10319_o ? 1'b1 : n10316_o;
  /* ppc_fx_insns.vhdl:758:22  */
  assign n10322_o = a_in[7:0];
  /* ppc_fx_insns.vhdl:758:39  */
  assign n10323_o = b_in[63:56];
  /* ppc_fx_insns.vhdl:758:35  */
  assign n10324_o = n10322_o == n10323_o;
  /* ppc_fx_insns.vhdl:758:17  */
  assign n10326_o = n10324_o ? 1'b1 : n10321_o;
  /* ppc_fx_insns.vhdl:762:24  */
  assign n10328_o = {1'b0, n10326_o};
  /* ppc_fx_insns.vhdl:762:32  */
  assign n10330_o = {n10328_o, 2'b00};
  /* execute1.vhdl:693:13  */
  assign n10332_o = n10226_o == 3'b010;
  /* execute1.vhdl:696:32  */
  assign n10333_o = current[344];
  /* execute1.vhdl:699:36  */
  assign n10342_o = 3'b111 - n10224_o;
  /* execute1.vhdl:700:40  */
  assign n10346_o = n9139_o[374:343];
  /* insn_helpers.vhdl:161:23  */
  assign n10351_o = n10346_o[25:21];
  /* execute1.vhdl:701:40  */
  assign n10353_o = n9139_o[374:343];
  /* insn_helpers.vhdl:156:23  */
  assign n10358_o = n10353_o[20:16];
  /* execute1.vhdl:702:40  */
  assign n10360_o = n9139_o[374:343];
  /* insn_helpers.vhdl:151:23  */
  assign n10365_o = n10360_o[15:11];
  /* execute1.vhdl:703:56  */
  assign n10366_o = n10351_o[1:0];
  /* execute1.vhdl:703:34  */
  assign n10367_o = {29'b0, n10366_o};  //  uext
  /* execute1.vhdl:703:32  */
  assign n10368_o = {1'b0, n10367_o};  //  uext
  /* execute1.vhdl:703:32  */
  assign n10370_o = 32'b00000000000000000000000000000011 - n10368_o;
  /* execute1.vhdl:703:21  */
  assign n10371_o = n10370_o[1:0];  // trunc
  /* execute1.vhdl:704:35  */
  assign n10372_o = {26'b0, n10358_o};  //  uext
  /* execute1.vhdl:704:33  */
  assign n10373_o = {1'b0, n10372_o};  //  uext
  /* execute1.vhdl:704:33  */
  assign n10375_o = 32'b00000000000000000000000000011111 - n10373_o;
  /* execute1.vhdl:704:21  */
  assign n10376_o = n10375_o[4:0];  // trunc
  /* execute1.vhdl:705:35  */
  assign n10377_o = {26'b0, n10365_o};  //  uext
  /* execute1.vhdl:705:33  */
  assign n10378_o = {1'b0, n10377_o};  //  uext
  /* execute1.vhdl:705:33  */
  assign n10380_o = 32'b00000000000000000000000000011111 - n10378_o;
  /* execute1.vhdl:705:21  */
  assign n10381_o = n10380_o[4:0];  // trunc
  /* execute1.vhdl:708:49  */
  assign n10386_o = {n12791_o, n12845_o};
  /* execute1.vhdl:709:47  */
  assign n10387_o = {29'b0, n10386_o};  //  uext
  /* execute1.vhdl:709:45  */
  assign n10388_o = {1'b0, n10387_o};  //  uext
  /* execute1.vhdl:709:45  */
  assign n10390_o = 32'b00000000000000000000000000000110 + n10388_o;
  /* execute1.vhdl:709:45  */
  assign n10391_o = n10390_o[4:0];  // trunc
  /* execute1.vhdl:711:30  */
  assign n10394_o = {30'b0, n10371_o};  //  uext
  /* execute1.vhdl:711:30  */
  assign n10396_o = 32'b00000000000000000000000000000000 == n10394_o;
  assign n10397_o = n12737_o[0];
  /* execute1.vhdl:711:25  */
  assign n10398_o = n10396_o ? n12899_o : n10397_o;
  /* execute1.vhdl:711:30  */
  assign n10400_o = {30'b0, n10371_o};  //  uext
  /* execute1.vhdl:711:30  */
  assign n10402_o = 32'b00000000000000000000000000000001 == n10400_o;
  assign n10403_o = n12737_o[1];
  /* execute1.vhdl:711:25  */
  assign n10404_o = n10402_o ? n12899_o : n10403_o;
  /* execute1.vhdl:711:30  */
  assign n10406_o = {30'b0, n10371_o};  //  uext
  /* execute1.vhdl:711:30  */
  assign n10408_o = 32'b00000000000000000000000000000010 == n10406_o;
  assign n10409_o = n12737_o[2];
  /* execute1.vhdl:711:25  */
  assign n10410_o = n10408_o ? n12899_o : n10409_o;
  assign n10411_o = n12737_o[3];
  /* execute1.vhdl:711:30  */
  assign n10412_o = {30'b0, n10371_o};  //  uext
  /* execute1.vhdl:711:30  */
  assign n10414_o = 32'b00000000000000000000000000000011 == n10412_o;
  /* execute1.vhdl:711:25  */
  assign n10415_o = n10414_o ? n12899_o : n10411_o;
  /* execute1.vhdl:717:42  */
  assign n10417_o = n9139_o[374:343];
  /* insn_helpers.vhdl:141:23  */
  assign n10422_o = n10417_o[20:18];
  /* execute1.vhdl:720:36  */
  assign n10432_o = 3'b111 - n10422_o;
  assign n10435_o = {n10415_o, n10410_o, n10404_o, n10398_o};
  /* execute1.vhdl:696:17  */
  assign n10436_o = n10333_o ? n10435_o : n12913_o;
  /* execute1.vhdl:695:13  */
  assign n10449_o = n10226_o == 3'b011;
  /* execute1.vhdl:724:35  */
  assign n10450_o = xerc_in[2];
  /* execute1.vhdl:724:48  */
  assign n10451_o = xerc_in[3];
  /* execute1.vhdl:724:38  */
  assign n10452_o = {n10450_o, n10451_o};
  /* execute1.vhdl:724:63  */
  assign n10453_o = xerc_in[0];
  /* execute1.vhdl:724:53  */
  assign n10454_o = {n10452_o, n10453_o};
  /* execute1.vhdl:724:76  */
  assign n10455_o = xerc_in[1];
  /* execute1.vhdl:724:66  */
  assign n10456_o = {n10454_o, n10455_o};
  /* execute1.vhdl:722:13  */
  assign n10458_o = n10226_o == 3'b100;
  assign n10459_o = {n10458_o, n10449_o, n10332_o, n10277_o, n10238_o};
  /* execute1.vhdl:683:9  */
  always @*
    case (n10459_o)
      5'b10000: n10461_o = n10456_o;
      5'b01000: n10461_o = n10436_o;
      5'b00100: n10461_o = n10330_o;
      5'b00010: n10461_o = n10275_o;
      5'b00001: n10461_o = n10236_o;
      default: n10461_o = 4'b0000;
    endcase
  /* execute1.vhdl:727:20  */
  assign n10474_o = current[9:4];
  /* execute1.vhdl:727:30  */
  assign n10476_o = n10474_o == 6'b100110;
  /* execute1.vhdl:728:25  */
  assign n10477_o = n9139_o[363];
  /* execute1.vhdl:728:30  */
  assign n10478_o = ~n10477_o;
  /* execute1.vhdl:730:48  */
  assign n10480_o = n9139_o[374:343];
  /* insn_helpers.vhdl:166:23  */
  assign n10485_o = n10480_o[19:12];
  /* execute1.vhdl:733:51  */
  assign n10488_o = n9139_o[374:343];
  /* insn_helpers.vhdl:166:23  */
  assign n10493_o = n10488_o[19:12];
  /* crhelpers.vhdl:23:19  */
  assign n10498_o = n10493_o[7];
  /* crhelpers.vhdl:23:13  */
  assign n10502_o = n10498_o ? 1'b0 : 1'b1;
  /* crhelpers.vhdl:23:13  */
  assign n10506_o = n10498_o ? 1'b0 : 1'b1;
  /* crhelpers.vhdl:23:13  */
  assign n10508_o = n10498_o ? 3'b000 : 3'bX;
  /* crhelpers.vhdl:23:19  */
  assign n10509_o = n10493_o[6];
  /* crhelpers.vhdl:23:13  */
  assign n10512_o = n10519_o ? 1'b0 : n10502_o;
  /* crhelpers.vhdl:23:13  */
  assign n10514_o = n10520_o ? 1'b0 : n10506_o;
  /* crhelpers.vhdl:23:13  */
  assign n10515_o = n10521_o ? 3'b001 : n10508_o;
  /* crhelpers.vhdl:23:13  */
  assign n10516_o = n10509_o & n10502_o;
  /* crhelpers.vhdl:23:13  */
  assign n10517_o = n10509_o & n10502_o;
  /* crhelpers.vhdl:23:13  */
  assign n10518_o = n10509_o & n10502_o;
  /* crhelpers.vhdl:23:13  */
  assign n10519_o = n10502_o & n10516_o;
  /* crhelpers.vhdl:23:13  */
  assign n10520_o = n10502_o & n10517_o;
  /* crhelpers.vhdl:23:13  */
  assign n10521_o = n10502_o & n10518_o;
  /* crhelpers.vhdl:23:19  */
  assign n10522_o = n10493_o[5];
  /* crhelpers.vhdl:23:13  */
  assign n10525_o = n10532_o ? 1'b0 : n10512_o;
  /* crhelpers.vhdl:23:13  */
  assign n10527_o = n10533_o ? 1'b0 : n10514_o;
  /* crhelpers.vhdl:23:13  */
  assign n10528_o = n10534_o ? 3'b010 : n10515_o;
  /* crhelpers.vhdl:23:13  */
  assign n10529_o = n10522_o & n10512_o;
  /* crhelpers.vhdl:23:13  */
  assign n10530_o = n10522_o & n10512_o;
  /* crhelpers.vhdl:23:13  */
  assign n10531_o = n10522_o & n10512_o;
  /* crhelpers.vhdl:23:13  */
  assign n10532_o = n10512_o & n10529_o;
  /* crhelpers.vhdl:23:13  */
  assign n10533_o = n10512_o & n10530_o;
  /* crhelpers.vhdl:23:13  */
  assign n10534_o = n10512_o & n10531_o;
  /* crhelpers.vhdl:23:19  */
  assign n10535_o = n10493_o[4];
  /* crhelpers.vhdl:23:13  */
  assign n10538_o = n10545_o ? 1'b0 : n10525_o;
  /* crhelpers.vhdl:23:13  */
  assign n10540_o = n10546_o ? 1'b0 : n10527_o;
  /* crhelpers.vhdl:23:13  */
  assign n10541_o = n10547_o ? 3'b011 : n10528_o;
  /* crhelpers.vhdl:23:13  */
  assign n10542_o = n10535_o & n10525_o;
  /* crhelpers.vhdl:23:13  */
  assign n10543_o = n10535_o & n10525_o;
  /* crhelpers.vhdl:23:13  */
  assign n10544_o = n10535_o & n10525_o;
  /* crhelpers.vhdl:23:13  */
  assign n10545_o = n10525_o & n10542_o;
  /* crhelpers.vhdl:23:13  */
  assign n10546_o = n10525_o & n10543_o;
  /* crhelpers.vhdl:23:13  */
  assign n10547_o = n10525_o & n10544_o;
  /* crhelpers.vhdl:23:19  */
  assign n10548_o = n10493_o[3];
  /* crhelpers.vhdl:23:13  */
  assign n10551_o = n10558_o ? 1'b0 : n10538_o;
  /* crhelpers.vhdl:23:13  */
  assign n10553_o = n10559_o ? 1'b0 : n10540_o;
  /* crhelpers.vhdl:23:13  */
  assign n10554_o = n10560_o ? 3'b100 : n10541_o;
  /* crhelpers.vhdl:23:13  */
  assign n10555_o = n10548_o & n10538_o;
  /* crhelpers.vhdl:23:13  */
  assign n10556_o = n10548_o & n10538_o;
  /* crhelpers.vhdl:23:13  */
  assign n10557_o = n10548_o & n10538_o;
  /* crhelpers.vhdl:23:13  */
  assign n10558_o = n10538_o & n10555_o;
  /* crhelpers.vhdl:23:13  */
  assign n10559_o = n10538_o & n10556_o;
  /* crhelpers.vhdl:23:13  */
  assign n10560_o = n10538_o & n10557_o;
  /* crhelpers.vhdl:23:19  */
  assign n10561_o = n10493_o[2];
  /* crhelpers.vhdl:23:13  */
  assign n10564_o = n10571_o ? 1'b0 : n10551_o;
  /* crhelpers.vhdl:23:13  */
  assign n10566_o = n10572_o ? 1'b0 : n10553_o;
  /* crhelpers.vhdl:23:13  */
  assign n10567_o = n10573_o ? 3'b101 : n10554_o;
  /* crhelpers.vhdl:23:13  */
  assign n10568_o = n10561_o & n10551_o;
  /* crhelpers.vhdl:23:13  */
  assign n10569_o = n10561_o & n10551_o;
  /* crhelpers.vhdl:23:13  */
  assign n10570_o = n10561_o & n10551_o;
  /* crhelpers.vhdl:23:13  */
  assign n10571_o = n10551_o & n10568_o;
  /* crhelpers.vhdl:23:13  */
  assign n10572_o = n10551_o & n10569_o;
  /* crhelpers.vhdl:23:13  */
  assign n10573_o = n10551_o & n10570_o;
  /* crhelpers.vhdl:23:19  */
  assign n10574_o = n10493_o[1];
  /* crhelpers.vhdl:23:13  */
  assign n10577_o = n10584_o ? 1'b0 : n10564_o;
  /* crhelpers.vhdl:23:13  */
  assign n10579_o = n10585_o ? 1'b0 : n10566_o;
  /* crhelpers.vhdl:23:13  */
  assign n10580_o = n10586_o ? 3'b110 : n10567_o;
  /* crhelpers.vhdl:23:13  */
  assign n10581_o = n10574_o & n10564_o;
  /* crhelpers.vhdl:23:13  */
  assign n10582_o = n10574_o & n10564_o;
  /* crhelpers.vhdl:23:13  */
  assign n10583_o = n10574_o & n10564_o;
  /* crhelpers.vhdl:23:13  */
  assign n10584_o = n10564_o & n10581_o;
  /* crhelpers.vhdl:23:13  */
  assign n10585_o = n10564_o & n10582_o;
  /* crhelpers.vhdl:23:13  */
  assign n10586_o = n10564_o & n10583_o;
  /* crhelpers.vhdl:23:19  */
  assign n10587_o = n10493_o[0];
  /* crhelpers.vhdl:23:13  */
  assign n10592_o = n10598_o ? 1'b0 : n10579_o;
  /* crhelpers.vhdl:23:13  */
  assign n10593_o = n10599_o ? 3'b111 : n10580_o;
  /* crhelpers.vhdl:23:13  */
  assign n10595_o = n10587_o & n10577_o;
  /* crhelpers.vhdl:23:13  */
  assign n10596_o = n10587_o & n10577_o;
  /* crhelpers.vhdl:23:13  */
  assign n10598_o = n10577_o & n10595_o;
  /* crhelpers.vhdl:23:13  */
  assign n10599_o = n10577_o & n10596_o;
  /* crhelpers.vhdl:30:9  */
  assign n10605_o = n10592_o ? 3'b111 : n10593_o;
  /* crhelpers.vhdl:36:13  */
  assign n10613_o = n10605_o == 3'b000;
  /* crhelpers.vhdl:38:13  */
  assign n10616_o = n10605_o == 3'b001;
  /* crhelpers.vhdl:40:13  */
  assign n10619_o = n10605_o == 3'b010;
  /* crhelpers.vhdl:42:13  */
  assign n10622_o = n10605_o == 3'b011;
  /* crhelpers.vhdl:44:13  */
  assign n10625_o = n10605_o == 3'b100;
  /* crhelpers.vhdl:46:13  */
  assign n10628_o = n10605_o == 3'b101;
  /* crhelpers.vhdl:48:13  */
  assign n10631_o = n10605_o == 3'b110;
  /* crhelpers.vhdl:50:13  */
  assign n10634_o = n10605_o == 3'b111;
  assign n10636_o = {n10634_o, n10631_o, n10628_o, n10625_o, n10622_o, n10619_o, n10616_o, n10613_o};
  /* crhelpers.vhdl:35:9  */
  always @*
    case (n10636_o)
      8'b10000000: n10637_o = 8'b00000001;
      8'b01000000: n10637_o = 8'b00000010;
      8'b00100000: n10637_o = 8'b00000100;
      8'b00010000: n10637_o = 8'b00001000;
      8'b00001000: n10637_o = 8'b00010000;
      8'b00000100: n10637_o = 8'b00100000;
      8'b00000010: n10637_o = 8'b01000000;
      8'b00000001: n10637_o = 8'b10000000;
      default: n10637_o = 8'b00000000;
    endcase
  /* execute1.vhdl:728:13  */
  assign n10638_o = n10478_o ? n10485_o : n10637_o;
  /* execute1.vhdl:736:34  */
  assign n10640_o = c_in[31:0];
  /* crhelpers.vhdl:36:13  */
  assign n10648_o = n10224_o == 3'b000;
  /* crhelpers.vhdl:38:13  */
  assign n10651_o = n10224_o == 3'b001;
  /* crhelpers.vhdl:40:13  */
  assign n10654_o = n10224_o == 3'b010;
  /* crhelpers.vhdl:42:13  */
  assign n10657_o = n10224_o == 3'b011;
  /* crhelpers.vhdl:44:13  */
  assign n10660_o = n10224_o == 3'b100;
  /* crhelpers.vhdl:46:13  */
  assign n10663_o = n10224_o == 3'b101;
  /* crhelpers.vhdl:48:13  */
  assign n10666_o = n10224_o == 3'b110;
  /* crhelpers.vhdl:50:13  */
  assign n10669_o = n10224_o == 3'b111;
  assign n10671_o = {n10669_o, n10666_o, n10663_o, n10660_o, n10657_o, n10654_o, n10651_o, n10648_o};
  /* crhelpers.vhdl:35:9  */
  always @*
    case (n10671_o)
      8'b10000000: n10672_o = 8'b00000001;
      8'b01000000: n10672_o = 8'b00000010;
      8'b00100000: n10672_o = 8'b00000100;
      8'b00010000: n10672_o = 8'b00001000;
      8'b00001000: n10672_o = 8'b00010000;
      8'b00000100: n10672_o = 8'b00100000;
      8'b00000010: n10672_o = 8'b01000000;
      8'b00000001: n10672_o = 8'b10000000;
      default: n10672_o = 8'b00000000;
    endcase
  /* execute1.vhdl:739:37  */
  assign n10673_o = {n10461_o, n10461_o};
  /* execute1.vhdl:739:46  */
  assign n10674_o = {n10673_o, n10461_o};
  /* execute1.vhdl:739:55  */
  assign n10675_o = {n10674_o, n10461_o};
  /* execute1.vhdl:739:64  */
  assign n10676_o = {n10675_o, n10461_o};
  /* execute1.vhdl:740:37  */
  assign n10677_o = {n10676_o, n10461_o};
  /* execute1.vhdl:740:46  */
  assign n10678_o = {n10677_o, n10461_o};
  /* execute1.vhdl:740:55  */
  assign n10679_o = {n10678_o, n10461_o};
  /* execute1.vhdl:727:9  */
  assign n10680_o = n10476_o ? n10638_o : n10672_o;
  /* execute1.vhdl:727:9  */
  assign n10681_o = n10476_o ? n10640_o : n10679_o;
  /* execute1.vhdl:770:35  */
  assign n10706_o = ctrl[133];
  /* execute1.vhdl:770:58  */
  assign n10707_o = ctrl[142];
  /* execute1.vhdl:770:46  */
  assign n10708_o = ~n10707_o;
  /* execute1.vhdl:770:44  */
  assign n10709_o = {n10706_o, n10708_o};
  /* execute1.vhdl:771:39  */
  assign n10710_o = ctrl[128];
  /* execute1.vhdl:771:27  */
  assign n10711_o = ~n10710_o;
  /* execute1.vhdl:770:67  */
  assign n10712_o = {n10709_o, n10711_o};
  /* execute1.vhdl:771:62  */
  assign n10713_o = ctrl[191];
  /* execute1.vhdl:771:50  */
  assign n10714_o = ~n10713_o;
  /* execute1.vhdl:771:48  */
  assign n10715_o = {n10712_o, n10714_o};
  assign n10737_o = r[798:767];
  /* execute1.vhdl:789:38  */
  assign n10740_o = ctrl[16];
  /* execute1.vhdl:790:38  */
  assign n10741_o = ctrl[12];
  /* execute1.vhdl:791:38  */
  assign n10742_o = ctrl[8];
  /* execute1.vhdl:792:38  */
  assign n10743_o = ctrl[0];
  /* execute1.vhdl:793:37  */
  assign n10744_o = ctrl[130];
  /* execute1.vhdl:794:36  */
  assign n10745_o = ctrl[142];
  /* execute1.vhdl:801:56  */
  assign n10746_o = ctrl[63:0];
  /* execute1.vhdl:801:60  */
  assign n10748_o = n10746_o + 64'b0000000000000000000000000000000000000000000000000000000000000001;
  /* execute1.vhdl:802:57  */
  assign n10750_o = ctrl[127:64];
  /* execute1.vhdl:802:62  */
  assign n10752_o = n10750_o - 64'b0000000000000000000000000000000000000000000000000000000000000001;
  assign n10753_o = ctrl[255:128];
  /* execute1.vhdl:804:30  */
  assign n10754_o = ctrl[143];
  /* execute1.vhdl:804:53  */
  assign n10755_o = pmu_to_x[64];
  /* execute1.vhdl:804:69  */
  assign n10756_o = ctrl[127];
  /* execute1.vhdl:804:58  */
  assign n10757_o = n10755_o | n10756_o;
  /* execute1.vhdl:804:74  */
  assign n10758_o = n10757_o | ext_irq_in;
  /* execute1.vhdl:804:39  */
  assign n10759_o = n10754_o & n10758_o;
  assign n10764_o = r[745:354];
  /* execute1.vhdl:811:53  */
  assign n10765_o = n9139_o[73:10];
  /* execute1.vhdl:811:58  */
  assign n10767_o = n10765_o + 64'b0000000000000000000000000000000000000000000000000000000000000100;
  /* execute1.vhdl:814:38  */
  assign n10769_o = n9139_o[9:4];
  /* execute1.vhdl:814:48  */
  assign n10771_o = n10769_o == 6'b110110;
  /* execute1.vhdl:814:28  */
  assign n10772_o = n10771_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:815:41  */
  assign n10775_o = n9139_o[9:4];
  /* execute1.vhdl:815:51  */
  assign n10777_o = n10775_o == 6'b110000;
  /* execute1.vhdl:815:68  */
  assign n10778_o = n9139_o[9:4];
  /* execute1.vhdl:815:78  */
  assign n10780_o = n10778_o == 6'b110001;
  /* execute1.vhdl:815:60  */
  assign n10781_o = n10777_o | n10780_o;
  /* execute1.vhdl:815:31  */
  assign n10782_o = n10781_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:816:42  */
  assign n10785_o = n9139_o[9:4];
  /* execute1.vhdl:816:52  */
  assign n10787_o = n10785_o == 6'b110000;
  /* execute1.vhdl:816:69  */
  assign n10788_o = n9139_o[9:4];
  /* execute1.vhdl:816:79  */
  assign n10790_o = n10788_o == 6'b110010;
  /* execute1.vhdl:816:61  */
  assign n10791_o = n10787_o | n10790_o;
  /* execute1.vhdl:816:32  */
  assign n10792_o = n10791_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:817:39  */
  assign n10795_o = n9139_o[9:4];
  /* execute1.vhdl:817:49  */
  assign n10797_o = n10795_o == 6'b011000;
  /* execute1.vhdl:817:29  */
  assign n10798_o = n10797_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:819:36  */
  assign n10801_o = n9139_o[9:4];
  /* execute1.vhdl:819:46  */
  assign n10803_o = n10801_o == 6'b101101;
  /* execute1.vhdl:819:26  */
  assign n10804_o = n10803_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:822:14  */
  assign n10806_o = r[748];
  /* execute1.vhdl:824:31  */
  assign n10809_o = r[353:0];
  /* execute1.vhdl:824:33  */
  assign n10810_o = n10809_o[137:126];
  assign n10811_o = n10704_o[137:126];
  /* execute1.vhdl:822:9  */
  assign n10812_o = n10806_o ? n10810_o : n10811_o;
  assign n10815_o = n10704_o[138];
  assign n10816_o = n10704_o[125];
  assign n10817_o = n10704_o[353:290];
  /* execute1.vhdl:827:34  */
  assign n10819_o = n9139_o[73:10];
  /* execute1.vhdl:829:31  */
  assign n10820_o = r[353:0];
  /* execute1.vhdl:829:33  */
  assign n10821_o = n10820_o[206:143];
  /* execute1.vhdl:826:9  */
  assign n10822_o = valid_in ? n10819_o : n10821_o;
  assign n10823_o = n10704_o[273:207];
  /* execute1.vhdl:832:39  */
  assign n10824_o = ctrl[191];
  /* execute1.vhdl:832:27  */
  assign n10825_o = ~n10824_o;
  assign n10826_o = n10704_o[119:6];
  /* execute1.vhdl:833:34  */
  assign n10828_o = current[76:74];
  assign n10829_o = n10704_o[4];
  assign n10830_o = n10704_o[0];
  /* execute1.vhdl:835:42  */
  assign n10831_o = ctrl[138];
  /* execute1.vhdl:835:30  */
  assign n10832_o = valid_in & n10831_o;
  /* execute1.vhdl:838:31  */
  assign n10833_o = n9139_o[9:4];
  /* execute1.vhdl:836:9  */
  assign n10834_o = valid_in ? n9139_o : n10764_o;
  assign n10835_o = r[756:751];
  /* execute1.vhdl:836:9  */
  assign n10836_o = valid_in ? n10833_o : n10835_o;
  assign n10837_o = r[757];
  /* execute1.vhdl:843:24  */
  assign n10839_o = r[748];
  /* execute1.vhdl:844:36  */
  assign n10840_o = n9139_o[391];
  /* execute1.vhdl:844:43  */
  assign n10841_o = ~n10840_o;
  /* execute1.vhdl:844:27  */
  assign n10842_o = valid_in & n10841_o;
  /* execute1.vhdl:844:55  */
  assign n10843_o = r[748];
  /* execute1.vhdl:844:68  */
  assign n10844_o = ~n10843_o;
  /* execute1.vhdl:844:49  */
  assign n10845_o = n10842_o & n10844_o;
  /* execute1.vhdl:845:30  */
  assign n10846_o = r[749];
  /* execute1.vhdl:845:24  */
  assign n10848_o = 1'b1 & n10846_o;
  /* execute1.vhdl:852:21  */
  assign n10852_o = r[750];
  /* execute1.vhdl:858:22  */
  assign n10855_o = r[756:751];
  /* execute1.vhdl:858:30  */
  assign n10857_o = n10855_o == 6'b011111;
  /* execute1.vhdl:858:45  */
  assign n10858_o = r[756:751];
  /* execute1.vhdl:858:53  */
  assign n10860_o = n10858_o == 6'b011011;
  /* execute1.vhdl:858:40  */
  assign n10861_o = n10857_o | n10860_o;
  /* execute1.vhdl:858:68  */
  assign n10862_o = r[756:751];
  /* execute1.vhdl:858:76  */
  assign n10864_o = n10862_o == 6'b011100;
  /* execute1.vhdl:858:63  */
  assign n10865_o = n10861_o | n10864_o;
  /* execute1.vhdl:859:23  */
  assign n10866_o = r[756:751];
  /* execute1.vhdl:859:31  */
  assign n10868_o = n10866_o == 6'b010010;
  /* execute1.vhdl:858:86  */
  assign n10869_o = n10865_o | n10868_o;
  /* execute1.vhdl:859:46  */
  assign n10870_o = r[756:751];
  /* execute1.vhdl:859:54  */
  assign n10872_o = n10870_o == 6'b010001;
  /* execute1.vhdl:859:41  */
  assign n10873_o = n10869_o | n10872_o;
  /* execute1.vhdl:859:70  */
  assign n10874_o = r[756:751];
  /* execute1.vhdl:859:78  */
  assign n10876_o = n10874_o == 6'b010000;
  /* execute1.vhdl:859:65  */
  assign n10877_o = n10873_o | n10876_o;
  /* execute1.vhdl:861:25  */
  assign n10879_o = r[756:751];
  /* execute1.vhdl:861:33  */
  assign n10881_o = n10879_o == 6'b100000;
  /* execute1.vhdl:861:49  */
  assign n10882_o = r[756:751];
  /* execute1.vhdl:861:57  */
  assign n10884_o = n10882_o == 6'b010100;
  /* execute1.vhdl:861:44  */
  assign n10885_o = n10881_o | n10884_o;
  /* execute1.vhdl:861:72  */
  assign n10886_o = r[756:751];
  /* execute1.vhdl:861:80  */
  assign n10888_o = n10886_o == 6'b010011;
  /* execute1.vhdl:861:67  */
  assign n10889_o = n10885_o | n10888_o;
  assign n10891_o = r[285];
  assign n10892_o = n10704_o[285];
  /* execute1.vhdl:822:9  */
  assign n10893_o = n10806_o ? n10891_o : n10892_o;
  /* execute1.vhdl:861:17  */
  assign n10894_o = n10889_o ? 1'b1 : n10893_o;
  assign n10895_o = r[285];
  assign n10896_o = n10704_o[285];
  /* execute1.vhdl:822:9  */
  assign n10897_o = n10806_o ? n10895_o : n10896_o;
  /* execute1.vhdl:858:17  */
  assign n10898_o = n10877_o ? n10897_o : n10894_o;
  assign n10899_o = r[286];
  assign n10900_o = n10704_o[286];
  /* execute1.vhdl:822:9  */
  assign n10901_o = n10806_o ? n10899_o : n10900_o;
  /* execute1.vhdl:858:17  */
  assign n10902_o = n10877_o ? 1'b1 : n10901_o;
  /* execute1.vhdl:868:29  */
  assign n10903_o = pmu_to_x[64];
  /* execute1.vhdl:871:31  */
  assign n10905_o = ctrl[127];
  /* execute1.vhdl:874:17  */
  assign n10909_o = ext_irq_in ? 12'b010100000000 : n10812_o;
  /* execute1.vhdl:874:17  */
  assign n10910_o = ext_irq_in ? 1'b1 : 1'b0;
  /* execute1.vhdl:871:17  */
  assign n10911_o = n10905_o ? 12'b100100000000 : n10909_o;
  /* execute1.vhdl:871:17  */
  assign n10912_o = n10905_o ? 1'b0 : n10910_o;
  /* execute1.vhdl:868:17  */
  assign n10913_o = n10903_o ? 12'b111100000000 : n10911_o;
  /* execute1.vhdl:868:17  */
  assign n10914_o = n10903_o ? 1'b0 : n10912_o;
  /* execute1.vhdl:881:27  */
  assign n10915_o = ctrl[142];
  /* execute1.vhdl:881:71  */
  assign n10917_o = n9139_o[9:4];
  /* execute1.vhdl:881:87  */
  assign n10918_o = n9139_o[374:343];
  /* execute1.vhdl:166:25  */
  assign n10924_o = 6'b111101 - n10917_o;
  /* execute1.vhdl:166:29  */
  assign n10929_o = n12561_data == 1'b1;
  /* execute1.vhdl:168:18  */
  assign n10932_o = n10917_o == 6'b100100;
  /* execute1.vhdl:168:35  */
  assign n10934_o = n10917_o == 6'b101000;
  /* execute1.vhdl:168:29  */
  assign n10935_o = n10932_o | n10934_o;
  /* execute1.vhdl:169:24  */
  assign n10936_o = n10918_o[20];
  /* execute1.vhdl:168:9  */
  assign n10938_o = n10935_o ? n10936_o : 1'b0;
  /* execute1.vhdl:166:9  */
  assign n10939_o = n10929_o ? 1'b1 : n10938_o;
  /* execute1.vhdl:881:42  */
  assign n10940_o = n10915_o & n10939_o;
  /* execute1.vhdl:893:39  */
  assign n10943_o = ctrl[141];
  /* execute1.vhdl:893:48  */
  assign n10944_o = ~n10943_o;
  /* execute1.vhdl:893:27  */
  assign n10946_o = 1'b1 & n10944_o;
  /* execute1.vhdl:893:63  */
  assign n10947_o = n9139_o[3];
  /* execute1.vhdl:893:67  */
  assign n10949_o = n10947_o == 1'b1;
  /* execute1.vhdl:893:54  */
  assign n10950_o = n10946_o & n10949_o;
  /* execute1.vhdl:893:13  */
  assign n10952_o = n10950_o ? 12'b100000000000 : n10812_o;
  /* execute1.vhdl:893:13  */
  assign n10954_o = n10950_o ? 1'b1 : n10839_o;
  /* execute1.vhdl:881:13  */
  assign n10955_o = n10940_o ? 12'b011100000000 : n10952_o;
  assign n10956_o = r[276];
  assign n10957_o = n10704_o[276];
  /* execute1.vhdl:822:9  */
  assign n10958_o = n10806_o ? n10956_o : n10957_o;
  /* execute1.vhdl:881:13  */
  assign n10959_o = n10940_o ? 1'b1 : n10958_o;
  /* execute1.vhdl:881:13  */
  assign n10961_o = n10940_o ? 1'b1 : n10954_o;
  /* execute1.vhdl:865:13  */
  assign n10962_o = n10759_o ? n10913_o : n10955_o;
  assign n10963_o = r[276];
  assign n10964_o = n10704_o[276];
  /* execute1.vhdl:822:9  */
  assign n10965_o = n10806_o ? n10963_o : n10964_o;
  /* execute1.vhdl:865:13  */
  assign n10966_o = n10759_o ? n10965_o : n10959_o;
  /* execute1.vhdl:865:13  */
  assign n10967_o = n10759_o ? n10914_o : 1'b0;
  /* execute1.vhdl:865:13  */
  assign n10969_o = n10759_o ? 1'b1 : n10961_o;
  assign n10970_o = {n10902_o, n10898_o};
  /* execute1.vhdl:852:13  */
  assign n10971_o = n10852_o ? 12'b110100000000 : n10962_o;
  assign n10972_o = r[276];
  assign n10973_o = n10704_o[276];
  /* execute1.vhdl:822:9  */
  assign n10974_o = n10806_o ? n10972_o : n10973_o;
  /* execute1.vhdl:852:13  */
  assign n10975_o = n10852_o ? n10974_o : n10966_o;
  assign n10976_o = r[286:285];
  assign n10977_o = n10704_o[286:285];
  /* execute1.vhdl:822:9  */
  assign n10978_o = n10806_o ? n10976_o : n10977_o;
  /* execute1.vhdl:852:13  */
  assign n10979_o = n10852_o ? n10970_o : n10978_o;
  assign n10980_o = r[288];
  assign n10981_o = n10704_o[288];
  /* execute1.vhdl:822:9  */
  assign n10982_o = n10806_o ? n10980_o : n10981_o;
  /* execute1.vhdl:852:13  */
  assign n10983_o = n10852_o ? 1'b1 : n10982_o;
  /* execute1.vhdl:852:13  */
  assign n10984_o = n10852_o ? 1'b0 : n10967_o;
  /* execute1.vhdl:852:13  */
  assign n10986_o = n10852_o ? 1'b1 : n10969_o;
  /* execute1.vhdl:845:13  */
  assign n10987_o = n10848_o ? 12'b011100000000 : n10971_o;
  assign n10988_o = r[274];
  assign n10989_o = n10704_o[274];
  /* execute1.vhdl:822:9  */
  assign n10990_o = n10806_o ? n10988_o : n10989_o;
  /* execute1.vhdl:845:13  */
  assign n10991_o = n10848_o ? 1'b1 : n10990_o;
  assign n10992_o = r[276];
  assign n10993_o = n10704_o[276];
  /* execute1.vhdl:822:9  */
  assign n10994_o = n10806_o ? n10992_o : n10993_o;
  /* execute1.vhdl:845:13  */
  assign n10995_o = n10848_o ? n10994_o : n10975_o;
  assign n10996_o = r[278];
  assign n10997_o = n10704_o[278];
  /* execute1.vhdl:822:9  */
  assign n10998_o = n10806_o ? n10996_o : n10997_o;
  /* execute1.vhdl:845:13  */
  assign n10999_o = n10848_o ? 1'b1 : n10998_o;
  assign n11000_o = r[286:285];
  assign n11001_o = n10704_o[286:285];
  /* execute1.vhdl:822:9  */
  assign n11002_o = n10806_o ? n11000_o : n11001_o;
  /* execute1.vhdl:845:13  */
  assign n11003_o = n10848_o ? n11002_o : n10979_o;
  assign n11004_o = r[288];
  assign n11005_o = n10704_o[288];
  /* execute1.vhdl:822:9  */
  assign n11006_o = n10806_o ? n11004_o : n11005_o;
  /* execute1.vhdl:845:13  */
  assign n11007_o = n10848_o ? n11006_o : n10983_o;
  /* execute1.vhdl:845:13  */
  assign n11008_o = n10848_o ? 1'b0 : n10984_o;
  /* execute1.vhdl:845:13  */
  assign n11010_o = n10848_o ? 1'b1 : n10986_o;
  /* execute1.vhdl:844:9  */
  assign n11011_o = n10845_o ? n10987_o : n10812_o;
  assign n11012_o = r[274];
  assign n11013_o = n10704_o[274];
  /* execute1.vhdl:822:9  */
  assign n11014_o = n10806_o ? n11012_o : n11013_o;
  /* execute1.vhdl:844:9  */
  assign n11015_o = n10845_o ? n10991_o : n11014_o;
  assign n11016_o = r[276];
  assign n11017_o = n10704_o[276];
  /* execute1.vhdl:822:9  */
  assign n11018_o = n10806_o ? n11016_o : n11017_o;
  /* execute1.vhdl:844:9  */
  assign n11019_o = n10845_o ? n10995_o : n11018_o;
  assign n11020_o = r[278];
  assign n11021_o = n10704_o[278];
  /* execute1.vhdl:822:9  */
  assign n11022_o = n10806_o ? n11020_o : n11021_o;
  /* execute1.vhdl:844:9  */
  assign n11023_o = n10845_o ? n10999_o : n11022_o;
  assign n11024_o = r[286:285];
  assign n11025_o = n10704_o[286:285];
  /* execute1.vhdl:822:9  */
  assign n11026_o = n10806_o ? n11024_o : n11025_o;
  /* execute1.vhdl:844:9  */
  assign n11027_o = n10845_o ? n11003_o : n11026_o;
  assign n11028_o = r[288];
  assign n11029_o = n10704_o[288];
  /* execute1.vhdl:822:9  */
  assign n11030_o = n10806_o ? n11028_o : n11029_o;
  /* execute1.vhdl:844:9  */
  assign n11031_o = n10845_o ? n11007_o : n11030_o;
  /* execute1.vhdl:844:9  */
  assign n11032_o = n10845_o ? n11008_o : 1'b0;
  assign n11039_o = r[275];
  assign n11040_o = n10704_o[275];
  /* execute1.vhdl:822:9  */
  assign n11041_o = n10806_o ? n11039_o : n11040_o;
  assign n11045_o = r[277];
  assign n11046_o = n10704_o[277];
  /* execute1.vhdl:822:9  */
  assign n11047_o = n10806_o ? n11045_o : n11046_o;
  assign n11051_o = r[284:279];
  assign n11052_o = n10704_o[284:279];
  /* execute1.vhdl:822:9  */
  assign n11053_o = n10806_o ? n11051_o : n11052_o;
  assign n11054_o = r[289];
  assign n11055_o = n10704_o[289];
  /* execute1.vhdl:822:9  */
  assign n11056_o = n10806_o ? n11054_o : n11055_o;
  assign n11057_o = r[287];
  assign n11058_o = n10704_o[287];
  /* execute1.vhdl:822:9  */
  assign n11059_o = n10806_o ? n11057_o : n11058_o;
  /* execute1.vhdl:844:9  */
  assign n11060_o = n10845_o ? n11010_o : n10839_o;
  /* execute1.vhdl:900:37  */
  assign n11061_o = n9140_o[1];
  /* execute1.vhdl:900:28  */
  assign n11062_o = n11060_o & n11061_o;
  /* execute1.vhdl:900:9  */
  assign n11065_o = n11062_o ? 1'b1 : 1'b0;
  assign n11066_o = r[748];
  /* execute1.vhdl:900:9  */
  assign n11067_o = n11062_o ? 1'b1 : n11066_o;
  assign n11068_o = r[750:749];
  /* execute1.vhdl:906:17  */
  assign n11069_o = n9140_o[2];
  /* execute1.vhdl:906:9  */
  assign n11071_o = n11069_o ? 1'b0 : n11067_o;
  /* execute1.vhdl:910:39  */
  assign n11072_o = n9139_o[0];
  /* execute1.vhdl:910:53  */
  assign n11073_o = n9140_o[0];
  /* execute1.vhdl:910:45  */
  assign n11074_o = n11072_o | n11073_o;
  /* execute1.vhdl:910:66  */
  assign n11075_o = n9140_o[1];
  /* execute1.vhdl:910:58  */
  assign n11076_o = n11074_o | n11075_o;
  /* execute1.vhdl:910:83  */
  assign n11077_o = r[746];
  /* execute1.vhdl:910:78  */
  assign n11078_o = n11076_o | n11077_o;
  /* execute1.vhdl:910:97  */
  assign n11079_o = n9141_o[0];
  /* execute1.vhdl:910:88  */
  assign n11080_o = n11078_o | n11079_o;
  /* execute1.vhdl:910:29  */
  assign n11081_o = ~n11080_o;
  /* execute1.vhdl:911:42  */
  assign n11083_o = ~n11060_o;
  /* execute1.vhdl:911:38  */
  assign n11084_o = valid_in & n11083_o;
  /* execute1.vhdl:911:56  */
  assign n11086_o = n11084_o & 1'b1;
  /* execute1.vhdl:913:41  */
  assign n11087_o = ~n11060_o;
  /* execute1.vhdl:913:27  */
  assign n11088_o = valid_in & n11087_o;
  /* execute1.vhdl:913:47  */
  assign n11090_o = n11088_o & 1'b1;
  /* execute1.vhdl:913:74  */
  assign n11091_o = n9139_o[2:1];
  /* execute1.vhdl:913:79  */
  assign n11093_o = n11091_o == 2'b01;
  /* execute1.vhdl:913:65  */
  assign n11094_o = n11090_o & n11093_o;
  /* execute1.vhdl:916:31  */
  assign n11096_o = n9139_o[9:4];
  /* execute1.vhdl:918:13  */
  assign n11098_o = n11096_o == 6'b000000;
  /* execute1.vhdl:926:29  */
  assign n11099_o = n9139_o[344];
  /* execute1.vhdl:926:17  */
  assign n11101_o = n11099_o ? 12'b110000000000 : n11011_o;
  /* execute1.vhdl:926:17  */
  assign n11102_o = n11099_o ? next_nia : n10822_o;
  /* execute1.vhdl:926:17  */
  assign n11104_o = n11099_o ? 1'b1 : n11060_o;
  /* execute1.vhdl:926:17  */
  assign n11107_o = n11099_o ? 1'b0 : 1'b1;
  /* execute1.vhdl:922:13  */
  assign n11109_o = n11096_o == 6'b110011;
  /* execute1.vhdl:937:29  */
  assign n11110_o = n9139_o[353:344];
  /* execute1.vhdl:937:43  */
  assign n11112_o = n11110_o == 10'b0100000000;
  /* execute1.vhdl:937:17  */
  assign n11114_o = n11112_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:937:17  */
  assign n11117_o = n11112_o ? 1'b0 : 1'b1;
  /* execute1.vhdl:934:13  */
  assign n11119_o = n11096_o == 6'b000100;
  /* execute1.vhdl:943:13  */
  assign n11121_o = n11096_o == 6'b000001;
  /* execute1.vhdl:943:25  */
  assign n11123_o = n11096_o == 6'b010000;
  /* execute1.vhdl:943:25  */
  assign n11124_o = n11121_o | n11123_o;
  /* execute1.vhdl:943:35  */
  assign n11126_o = n11096_o == 6'b010001;
  /* execute1.vhdl:943:35  */
  assign n11127_o = n11124_o | n11126_o;
  /* execute1.vhdl:943:46  */
  assign n11129_o = n11096_o == 6'b010010;
  /* execute1.vhdl:943:46  */
  assign n11130_o = n11127_o | n11129_o;
  /* execute1.vhdl:943:56  */
  assign n11132_o = n11096_o == 6'b010011;
  /* execute1.vhdl:943:56  */
  assign n11133_o = n11130_o | n11132_o;
  /* execute1.vhdl:943:68  */
  assign n11135_o = n11096_o == 6'b011100;
  /* execute1.vhdl:943:68  */
  assign n11136_o = n11133_o | n11135_o;
  /* execute1.vhdl:946:25  */
  assign n11137_o = n9139_o[337];
  /* execute1.vhdl:947:29  */
  assign n11138_o = n9139_o[336:335];
  /* execute1.vhdl:947:41  */
  assign n11140_o = n11138_o != 2'b10;
  assign n11142_o = {n10737_o, 1'b0, 1'b0, n11032_o, n11086_o, n11081_o, 1'b0, 1'b0, 1'b0, 1'b0, n10837_o, n10836_o, n11068_o, n11071_o, 1'b0, n11065_o, n10834_o, n10817_o, n11056_o, n11031_o, n11059_o, n11027_o, n11053_o, n11023_o, n11047_o, n11019_o, n11041_o, n11015_o, n10823_o, n10822_o, n10715_o, n10815_o, n11011_o, n10816_o, xerc_in, n10826_o, n10825_o, n10829_o, n10828_o, 1'b1};
  assign n11146_o = n11142_o[119:0];
  assign n11147_o = n11142_o[353:122];
  assign n11148_o = {n11147_o, carry_32, carry_64, n11146_o};
  assign n11149_o = {carry_32, carry_64};
  assign n11150_o = n11148_o[121:0];
  assign n11151_o = xerc_in[1:0];
  assign n11152_o = {n11151_o, n10826_o, n10825_o, n10829_o, n10828_o, 1'b1};
  /* execute1.vhdl:947:21  */
  assign n11153_o = n11140_o ? n11150_o : n11152_o;
  assign n11154_o = n11148_o[123:122];
  /* execute1.vhdl:947:21  */
  assign n11155_o = n11140_o ? n11154_o : n11149_o;
  assign n11156_o = n11148_o[353:124];
  assign n11157_o = xerc_in[4];
  assign n11158_o = {n10817_o, n11056_o, n11031_o, n11059_o, n11027_o, n11053_o, n11023_o, n11047_o, n11019_o, n11041_o, n11015_o, n10823_o, n10822_o, n10715_o, n10815_o, n11011_o, n10816_o, n11157_o};
  /* execute1.vhdl:947:21  */
  assign n11159_o = n11140_o ? n11156_o : n11158_o;
  assign n11160_o = {n11159_o, n11155_o, n11153_o};
  assign n11161_o = {n10817_o, n11056_o, n11031_o, n11059_o, n11027_o, n11053_o, n11023_o, n11047_o, n11019_o, n11041_o, n11015_o, n10823_o, n10822_o, n10715_o, n10815_o, n11011_o, n10816_o, xerc_in, n10826_o, n10825_o, n10829_o, n10828_o, 1'b1};
  /* execute1.vhdl:946:17  */
  assign n11162_o = n11137_o ? n11160_o : n11161_o;
  /* execute1.vhdl:954:25  */
  assign n11163_o = n9139_o[331];
  assign n11165_o = {n10737_o, 1'b0, 1'b0, n11032_o, n11086_o, n11081_o, 1'b0, 1'b0, 1'b0, 1'b0, n10837_o, n10836_o, n11068_o, n11071_o, 1'b0, n11065_o, n10834_o, n11162_o};
  assign n11170_o = n11165_o[124];
  /* execute1.vhdl:189:9  */
  assign n11171_o = overflow_64 ? 1'b1 : n11170_o;
  assign n11172_o = n11165_o[121:0];
  assign n11173_o = n11165_o[353:125];
  assign n11174_o = {n11173_o, n11171_o, overflow_32, overflow_64, n11172_o};
  /* execute1.vhdl:954:17  */
  assign n11175_o = n11163_o ? n11174_o : n11162_o;
  /* execute1.vhdl:945:13  */
  assign n11177_o = n11096_o == 6'b000010;
  /* execute1.vhdl:957:13  */
  assign n11179_o = n11096_o == 6'b001001;
  /* execute1.vhdl:963:49  */
  assign n11183_o = n9139_o[374:343];
  /* insn_helpers.vhdl:206:23  */
  assign n11188_o = n11183_o[25:21];
  /* execute1.vhdl:963:32  */
  assign n11189_o = trapval & n11188_o;
  /* execute1.vhdl:963:20  */
  assign n11190_o = |(n11189_o);
  /* execute1.vhdl:963:17  */
  assign n11192_o = n11190_o ? 1'b1 : n11060_o;
  /* execute1.vhdl:958:13  */
  assign n11194_o = n11096_o == 6'b111001;
  /* execute1.vhdl:968:13  */
  assign n11196_o = n11096_o == 6'b111100;
  /* execute1.vhdl:969:13  */
  assign n11198_o = n11096_o == 6'b001100;
  /* execute1.vhdl:970:13  */
  assign n11200_o = n11096_o == 6'b001011;
  /* execute1.vhdl:971:13  */
  assign n11202_o = n11096_o == 6'b000011;
  /* execute1.vhdl:971:25  */
  assign n11204_o = n11096_o == 6'b101100;
  /* execute1.vhdl:971:25  */
  assign n11205_o = n11202_o | n11204_o;
  /* execute1.vhdl:971:33  */
  assign n11207_o = n11096_o == 6'b111010;
  /* execute1.vhdl:971:33  */
  assign n11208_o = n11205_o | n11207_o;
  /* execute1.vhdl:971:42  */
  assign n11210_o = n11096_o == 6'b101110;
  /* execute1.vhdl:971:42  */
  assign n11211_o = n11208_o | n11210_o;
  /* execute1.vhdl:971:52  */
  assign n11213_o = n11096_o == 6'b001010;
  /* execute1.vhdl:971:52  */
  assign n11214_o = n11211_o | n11213_o;
  /* execute1.vhdl:971:62  */
  assign n11216_o = n11096_o == 6'b010111;
  /* execute1.vhdl:971:62  */
  assign n11217_o = n11214_o | n11216_o;
  /* execute1.vhdl:971:72  */
  assign n11219_o = n11096_o == 6'b001000;
  /* execute1.vhdl:971:72  */
  assign n11220_o = n11217_o | n11219_o;
  /* execute1.vhdl:972:30  */
  assign n11222_o = n11096_o == 6'b111011;
  /* execute1.vhdl:972:30  */
  assign n11223_o = n11220_o | n11222_o;
  /* execute1.vhdl:978:36  */
  assign n11224_o = n9139_o[329];
  /* execute1.vhdl:979:28  */
  assign n11225_o = ctrl[137];
  /* execute1.vhdl:979:17  */
  assign n11227_o = n11225_o ? 1'b1 : n10832_o;
  /* execute1.vhdl:974:13  */
  assign n11230_o = n11096_o == 6'b000101;
  /* execute1.vhdl:990:36  */
  assign n11232_o = n9139_o[374:343];
  /* insn_helpers.vhdl:171:23  */
  assign n11237_o = n11232_o[25:21];
  /* execute1.vhdl:991:36  */
  assign n11239_o = n9139_o[374:343];
  /* insn_helpers.vhdl:176:23  */
  assign n11244_o = n11239_o[20:16];
  /* execute1.vhdl:992:25  */
  assign n11245_o = n9139_o[391];
  /* execute1.vhdl:992:32  */
  assign n11246_o = ~n11245_o;
  /* ppc_fx_insns.vhdl:825:28  */
  assign n11257_o = {26'b0, n11244_o};  //  uext
  /* ppc_fx_insns.vhdl:825:17  */
  assign n11258_o = {1'b0, n11257_o};  //  uext
  /* ppc_fx_insns.vhdl:827:46  */
  assign n11261_o = 32'b00000000000000000000000000011111 - n11258_o;
  /* ppc_fx_insns.vhdl:827:46  */
  assign n11262_o = n11261_o[4:0];  // trunc
  /* ppc_fx_insns.vhdl:827:60  */
  assign n11265_o = n11237_o[3];
  /* ppc_fx_insns.vhdl:827:56  */
  assign n11266_o = n12967_o == n11265_o;
  /* ppc_fx_insns.vhdl:827:36  */
  assign n11268_o = n11266_o ? 1'b1 : 1'b0;
  /* ppc_fx_insns.vhdl:829:46  */
  assign n11272_o = a_in != 64'b0000000000000000000000000000000000000000000000000000000000000001;
  /* ppc_fx_insns.vhdl:829:37  */
  assign n11274_o = n11272_o ? 1'b1 : 1'b0;
  /* ppc_fx_insns.vhdl:830:29  */
  assign n11277_o = n11237_o[2];
  /* ppc_fx_insns.vhdl:830:58  */
  assign n11278_o = n11237_o[1];
  /* ppc_fx_insns.vhdl:830:52  */
  assign n11279_o = n11274_o ^ n11278_o;
  /* ppc_fx_insns.vhdl:830:35  */
  assign n11280_o = n11277_o | n11279_o;
  /* ppc_fx_insns.vhdl:831:30  */
  assign n11282_o = n11237_o[4];
  /* ppc_fx_insns.vhdl:831:36  */
  assign n11283_o = n11282_o | n11268_o;
  /* ppc_fx_insns.vhdl:832:31  */
  assign n11285_o = n11280_o & n11283_o;
  /* execute1.vhdl:995:39  */
  assign n11286_o = r[757];
  /* execute1.vhdl:992:17  */
  assign n11287_o = n11246_o ? n11285_o : n11286_o;
  /* execute1.vhdl:999:36  */
  assign n11288_o = n9139_o[329];
  /* execute1.vhdl:1000:25  */
  assign n11289_o = n9139_o[390];
  /* execute1.vhdl:1000:32  */
  assign n11290_o = ~n11289_o;
  /* execute1.vhdl:1000:46  */
  assign n11291_o = n9139_o[391];
  /* execute1.vhdl:1000:38  */
  assign n11292_o = n11290_o | n11291_o;
  /* execute1.vhdl:1002:29  */
  assign n11293_o = n9139_o[9:4];
  /* execute1.vhdl:1002:39  */
  assign n11295_o = n11293_o == 6'b000110;
  /* execute1.vhdl:1002:21  */
  assign n11298_o = n11295_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:1005:32  */
  assign n11299_o = ctrl[137];
  /* execute1.vhdl:1000:17  */
  assign n11301_o = n11307_o ? 1'b1 : n10832_o;
  /* execute1.vhdl:1000:17  */
  assign n11304_o = n11292_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:1000:17  */
  assign n11306_o = n11292_o ? n11298_o : 1'b0;
  /* execute1.vhdl:1000:17  */
  assign n11307_o = n11292_o & n11299_o;
  /* execute1.vhdl:983:13  */
  assign n11309_o = n11096_o == 6'b000110;
  /* execute1.vhdl:983:24  */
  assign n11311_o = n11096_o == 6'b000111;
  /* execute1.vhdl:983:24  */
  assign n11312_o = n11309_o | n11311_o;
  /* execute1.vhdl:1011:40  */
  assign n11313_o = a_in[5];
  /* execute1.vhdl:1011:56  */
  assign n11314_o = a_in[14];
  /* execute1.vhdl:1011:49  */
  assign n11315_o = n11313_o | n11314_o;
  /* execute1.vhdl:1011:76  */
  assign n11316_o = a_in[14];
  /* execute1.vhdl:1011:68  */
  assign n11317_o = ~n11316_o;
  /* execute1.vhdl:1011:66  */
  assign n11318_o = {n11315_o, n11317_o};
  /* execute1.vhdl:1012:43  */
  assign n11319_o = a_in[0];
  /* execute1.vhdl:1012:35  */
  assign n11320_o = ~n11319_o;
  /* execute1.vhdl:1011:85  */
  assign n11321_o = {n11318_o, n11320_o};
  /* execute1.vhdl:1012:62  */
  assign n11322_o = a_in[63];
  /* execute1.vhdl:1012:54  */
  assign n11323_o = ~n11322_o;
  /* execute1.vhdl:1012:52  */
  assign n11324_o = {n11321_o, n11323_o};
  /* execute1.vhdl:1015:51  */
  assign n11325_o = a_in[63:31];
  /* execute1.vhdl:1016:51  */
  assign n11326_o = a_in[26:22];
  /* execute1.vhdl:1018:24  */
  assign n11328_o = a_in[14];
  assign n11332_o = {1'b1, 1'b1};
  assign n11333_o = a_in[5:4];
  /* execute1.vhdl:1018:17  */
  assign n11334_o = n11328_o ? n11332_o : n11333_o;
  assign n11335_o = a_in[15];
  /* execute1.vhdl:1018:17  */
  assign n11336_o = n11328_o ? 1'b1 : n11335_o;
  assign n11338_o = a_in[3:0];
  assign n11339_o = a_in[14:6];
  /* execute1.vhdl:1028:50  */
  assign n11340_o = n9141_o[1];
  /* execute1.vhdl:1029:49  */
  assign n11341_o = a_in[11];
  /* execute1.vhdl:1029:66  */
  assign n11342_o = a_in[8];
  /* execute1.vhdl:1029:59  */
  assign n11343_o = n11341_o | n11342_o;
  /* execute1.vhdl:1028:60  */
  assign n11344_o = n11340_o & n11343_o;
  /* execute1.vhdl:1010:13  */
  assign n11346_o = n11096_o == 6'b101111;
  /* execute1.vhdl:1033:13  */
  assign n11351_o = n11096_o == 6'b001101;
  /* execute1.vhdl:1033:26  */
  assign n11353_o = n11096_o == 6'b101101;
  /* execute1.vhdl:1033:26  */
  assign n11354_o = n11351_o | n11353_o;
  /* execute1.vhdl:1037:13  */
  assign n11356_o = n11096_o == 6'b011101;
  /* execute1.vhdl:1038:13  */
  assign n11358_o = n11096_o == 6'b001110;
  /* execute1.vhdl:1039:13  */
  assign n11360_o = n11096_o == 6'b100001;
  /* execute1.vhdl:1040:13  */
  assign n11362_o = n11096_o == 6'b001111;
  /* execute1.vhdl:1041:13  */
  assign n11364_o = n11096_o == 6'b100011;
  /* execute1.vhdl:1045:37  */
  assign n11366_o = n9139_o[91:85];
  /* common.vhdl:775:17  */
  assign n11371_o = n11366_o[5];
  /* execute1.vhdl:1047:44  */
  assign n11373_o = n9139_o[374:343];
  /* common.vhdl:708:40  */
  assign n11378_o = n11373_o[15:11];
  /* common.vhdl:708:61  */
  assign n11379_o = n11373_o[20:16];
  /* common.vhdl:708:55  */
  assign n11380_o = {n11378_o, n11379_o};
  /* execute1.vhdl:1047:50  */
  assign n11382_o = {22'b0, n11380_o};  //  uext
  /* execute1.vhdl:1047:50  */
  assign n11384_o = n11382_o == 32'b00000000000000000000000000000001;
  /* execute1.vhdl:1050:51  */
  assign n11386_o = xerc_in[4];
  /* execute1.vhdl:1051:51  */
  assign n11387_o = xerc_in[2];
  /* execute1.vhdl:1052:51  */
  assign n11388_o = xerc_in[0];
  /* execute1.vhdl:1054:51  */
  assign n11390_o = xerc_in[3];
  /* execute1.vhdl:1055:51  */
  assign n11391_o = xerc_in[1];
  assign n11392_o = {32'b00000000000000000000000000000000, n11386_o, n11387_o, n11388_o, 9'b000000000, n11390_o, n11391_o};
  assign n11393_o = a_in[63:18];
  /* execute1.vhdl:1047:21  */
  assign n11394_o = n11384_o ? n11392_o : n11393_o;
  assign n11395_o = a_in[17:0];
  /* execute1.vhdl:1059:46  */
  assign n11397_o = n9139_o[374:343];
  /* common.vhdl:708:40  */
  assign n11402_o = n11397_o[15:11];
  /* common.vhdl:708:61  */
  assign n11403_o = n11397_o[20:16];
  /* common.vhdl:708:55  */
  assign n11404_o = {n11402_o, n11403_o};
  /* execute1.vhdl:1061:41  */
  assign n11406_o = ctrl[63:0];
  /* execute1.vhdl:1060:21  */
  assign n11408_o = n11404_o == 10'b0100001100;
  /* execute1.vhdl:1064:57  */
  assign n11410_o = ctrl[63:32];
  /* execute1.vhdl:1062:21  */
  assign n11412_o = n11404_o == 10'b0100001101;
  /* execute1.vhdl:1066:41  */
  assign n11413_o = ctrl[127:64];
  /* execute1.vhdl:1065:21  */
  assign n11415_o = n11404_o == 10'b0000010110;
  /* execute1.vhdl:1068:41  */
  assign n11416_o = ctrl[255:192];
  /* execute1.vhdl:1067:21  */
  assign n11418_o = n11404_o == 10'b0000011100;
  /* execute1.vhdl:1069:21  */
  assign n11422_o = n11404_o == 10'b0100011111;
  /* execute1.vhdl:1073:52  */
  assign n11423_o = r[798:767];
  /* execute1.vhdl:1073:48  */
  assign n11424_o = {log_wr_addr, n11423_o};
  /* execute1.vhdl:1072:21  */
  assign n11426_o = n11404_o == 10'b1011010100;
  /* execute1.vhdl:1076:72  */
  assign n11427_o = r[798:767];
  /* execute1.vhdl:1076:86  */
  assign n11429_o = n11427_o + 32'b00000000000000000000000000000001;
  /* execute1.vhdl:1074:21  */
  assign n11431_o = n11404_o == 10'b1011010101;
  /* execute1.vhdl:1082:45  */
  assign n11433_o = pmu_to_x[63:0];
  /* execute1.vhdl:1077:21  */
  assign n11435_o = n11404_o == 10'b1100000011;
  /* execute1.vhdl:1077:36  */
  assign n11437_o = n11404_o == 10'b1100000100;
  /* execute1.vhdl:1077:36  */
  assign n11438_o = n11435_o | n11437_o;
  /* execute1.vhdl:1077:48  */
  assign n11440_o = n11404_o == 10'b1100000101;
  /* execute1.vhdl:1077:48  */
  assign n11441_o = n11438_o | n11440_o;
  /* execute1.vhdl:1077:60  */
  assign n11443_o = n11404_o == 10'b1100000110;
  /* execute1.vhdl:1077:60  */
  assign n11444_o = n11441_o | n11443_o;
  /* execute1.vhdl:1077:72  */
  assign n11446_o = n11404_o == 10'b1100000111;
  /* execute1.vhdl:1077:72  */
  assign n11447_o = n11444_o | n11446_o;
  /* execute1.vhdl:1077:84  */
  assign n11449_o = n11404_o == 10'b1100001000;
  /* execute1.vhdl:1077:84  */
  assign n11450_o = n11447_o | n11449_o;
  /* execute1.vhdl:1077:96  */
  assign n11452_o = n11404_o == 10'b1100001011;
  /* execute1.vhdl:1077:96  */
  assign n11453_o = n11450_o | n11452_o;
  /* execute1.vhdl:1078:36  */
  assign n11455_o = n11404_o == 10'b1100001110;
  /* execute1.vhdl:1078:36  */
  assign n11456_o = n11453_o | n11455_o;
  /* execute1.vhdl:1078:49  */
  assign n11458_o = n11404_o == 10'b1100000001;
  /* execute1.vhdl:1078:49  */
  assign n11459_o = n11456_o | n11458_o;
  /* execute1.vhdl:1078:62  */
  assign n11461_o = n11404_o == 10'b1100000010;
  /* execute1.vhdl:1078:62  */
  assign n11462_o = n11459_o | n11461_o;
  /* execute1.vhdl:1078:75  */
  assign n11464_o = n11404_o == 10'b1100000000;
  /* execute1.vhdl:1078:75  */
  assign n11465_o = n11462_o | n11464_o;
  /* execute1.vhdl:1078:87  */
  assign n11467_o = n11404_o == 10'b1100001100;
  /* execute1.vhdl:1078:87  */
  assign n11468_o = n11465_o | n11467_o;
  /* execute1.vhdl:1078:99  */
  assign n11470_o = n11404_o == 10'b1100001101;
  /* execute1.vhdl:1078:99  */
  assign n11471_o = n11468_o | n11470_o;
  /* execute1.vhdl:1078:111  */
  assign n11473_o = n11404_o == 10'b1100010011;
  /* execute1.vhdl:1078:111  */
  assign n11474_o = n11471_o | n11473_o;
  /* execute1.vhdl:1079:34  */
  assign n11476_o = n11404_o == 10'b1100010100;
  /* execute1.vhdl:1079:34  */
  assign n11477_o = n11474_o | n11476_o;
  /* execute1.vhdl:1079:45  */
  assign n11479_o = n11404_o == 10'b1100010101;
  /* execute1.vhdl:1079:45  */
  assign n11480_o = n11477_o | n11479_o;
  /* execute1.vhdl:1079:56  */
  assign n11482_o = n11404_o == 10'b1100010110;
  /* execute1.vhdl:1079:56  */
  assign n11483_o = n11480_o | n11482_o;
  /* execute1.vhdl:1079:67  */
  assign n11485_o = n11404_o == 10'b1100010111;
  /* execute1.vhdl:1079:67  */
  assign n11486_o = n11483_o | n11485_o;
  /* execute1.vhdl:1079:78  */
  assign n11488_o = n11404_o == 10'b1100011000;
  /* execute1.vhdl:1079:78  */
  assign n11489_o = n11486_o | n11488_o;
  /* execute1.vhdl:1079:89  */
  assign n11491_o = n11404_o == 10'b1100011011;
  /* execute1.vhdl:1079:89  */
  assign n11492_o = n11489_o | n11491_o;
  /* execute1.vhdl:1080:35  */
  assign n11494_o = n11404_o == 10'b1100011110;
  /* execute1.vhdl:1080:35  */
  assign n11495_o = n11492_o | n11494_o;
  /* execute1.vhdl:1080:47  */
  assign n11497_o = n11404_o == 10'b1100010001;
  /* execute1.vhdl:1080:47  */
  assign n11498_o = n11495_o | n11497_o;
  /* execute1.vhdl:1080:59  */
  assign n11500_o = n11404_o == 10'b1100010010;
  /* execute1.vhdl:1080:59  */
  assign n11501_o = n11498_o | n11500_o;
  /* execute1.vhdl:1080:71  */
  assign n11503_o = n11404_o == 10'b1100010000;
  /* execute1.vhdl:1080:71  */
  assign n11504_o = n11501_o | n11503_o;
  /* execute1.vhdl:1080:82  */
  assign n11506_o = n11404_o == 10'b1100011100;
  /* execute1.vhdl:1080:82  */
  assign n11507_o = n11504_o | n11506_o;
  /* execute1.vhdl:1080:93  */
  assign n11509_o = n11404_o == 10'b1100011101;
  /* execute1.vhdl:1080:93  */
  assign n11510_o = n11507_o | n11509_o;
  /* execute1.vhdl:1086:45  */
  assign n11512_o = n9139_o[91:85];
  /* common.vhdl:775:17  */
  assign n11517_o = n11512_o[5];
  /* execute1.vhdl:1086:56  */
  assign n11518_o = ~n11517_o;
  /* execute1.vhdl:1086:74  */
  assign n11519_o = ctrl[142];
  /* execute1.vhdl:1086:62  */
  assign n11520_o = n11518_o & n11519_o;
  /* execute1.vhdl:1086:25  */
  assign n11523_o = n11520_o ? 1'b1 : 1'b0;
  assign n11524_o = {n11510_o, n11431_o, n11426_o, n11422_o, n11418_o, n11415_o, n11412_o, n11408_o};
  /* execute1.vhdl:1059:21  */
  always @*
    case (n11524_o)
      8'b10000000: n11525_o = 1'b1;
      8'b01000000: n11525_o = 1'b0;
      8'b00100000: n11525_o = 1'b0;
      8'b00010000: n11525_o = 1'b0;
      8'b00001000: n11525_o = 1'b0;
      8'b00000100: n11525_o = 1'b0;
      8'b00000010: n11525_o = 1'b0;
      8'b00000001: n11525_o = 1'b0;
      default: n11525_o = 1'b0;
    endcase
  /* execute1.vhdl:1059:21  */
  always @*
    case (n11524_o)
      8'b10000000: n11526_o = n10737_o;
      8'b01000000: n11526_o = n11429_o;
      8'b00100000: n11526_o = n10737_o;
      8'b00010000: n11526_o = n10737_o;
      8'b00001000: n11526_o = n10737_o;
      8'b00000100: n11526_o = n10737_o;
      8'b00000010: n11526_o = n10737_o;
      8'b00000001: n11526_o = n10737_o;
      default: n11526_o = n10737_o;
    endcase
  /* execute1.vhdl:1059:21  */
  always @*
    case (n11524_o)
      8'b10000000: n11528_o = 1'b0;
      8'b01000000: n11528_o = 1'b0;
      8'b00100000: n11528_o = 1'b0;
      8'b00010000: n11528_o = 1'b0;
      8'b00001000: n11528_o = 1'b0;
      8'b00000100: n11528_o = 1'b0;
      8'b00000010: n11528_o = 1'b0;
      8'b00000001: n11528_o = 1'b0;
      default: n11528_o = n11523_o;
    endcase
  assign n11529_o = n11406_o[31:0];
  assign n11530_o = n11413_o[31:0];
  assign n11531_o = n11416_o[31:0];
  assign n11532_o = n11424_o[31:0];
  assign n11533_o = log_rd_data[31:0];
  assign n11534_o = n11433_o[31:0];
  assign n11535_o = c_in[31:0];
  /* execute1.vhdl:1059:21  */
  always @*
    case (n11524_o)
      8'b10000000: n11536_o = n11534_o;
      8'b01000000: n11536_o = n11533_o;
      8'b00100000: n11536_o = n11532_o;
      8'b00010000: n11536_o = 32'b00000000011000110000000100000001;
      8'b00001000: n11536_o = n11531_o;
      8'b00000100: n11536_o = n11530_o;
      8'b00000010: n11536_o = n11410_o;
      8'b00000001: n11536_o = n11529_o;
      default: n11536_o = n11535_o;
    endcase
  assign n11537_o = n11406_o[63:32];
  assign n11538_o = n11413_o[63:32];
  assign n11539_o = n11416_o[63:32];
  assign n11540_o = n11424_o[63:32];
  assign n11541_o = log_rd_data[63:32];
  assign n11542_o = n11433_o[63:32];
  assign n11543_o = c_in[63:32];
  /* execute1.vhdl:1059:21  */
  always @*
    case (n11524_o)
      8'b10000000: n11544_o = n11542_o;
      8'b01000000: n11544_o = n11541_o;
      8'b00100000: n11544_o = n11540_o;
      8'b00010000: n11544_o = 32'b00000000000000000000000000000000;
      8'b00001000: n11544_o = n11539_o;
      8'b00000100: n11544_o = n11538_o;
      8'b00000010: n11544_o = 32'b00000000000000000000000000000000;
      8'b00000001: n11544_o = n11537_o;
      default: n11544_o = n11543_o;
    endcase
  /* execute1.vhdl:1045:17  */
  assign n11546_o = n11371_o ? 1'b0 : n11525_o;
  /* execute1.vhdl:1045:17  */
  assign n11547_o = n11371_o ? n10737_o : n11526_o;
  /* execute1.vhdl:1045:17  */
  assign n11549_o = n11371_o ? 1'b0 : n11528_o;
  assign n11550_o = {n11544_o, n11536_o};
  assign n11551_o = {n11394_o, n11395_o};
  /* execute1.vhdl:1045:17  */
  assign n11552_o = n11371_o ? n11551_o : n11550_o;
  /* execute1.vhdl:1042:13  */
  assign n11554_o = n11096_o == 6'b100100;
  /* execute1.vhdl:1093:13  */
  assign n11556_o = n11096_o == 6'b100010;
  /* execute1.vhdl:1094:13  */
  assign n11558_o = n11096_o == 6'b100110;
  /* execute1.vhdl:1096:29  */
  assign n11559_o = n9139_o[359];
  /* execute1.vhdl:1098:49  */
  assign n11560_o = c_in[15];
  /* execute1.vhdl:1099:49  */
  assign n11561_o = c_in[1];
  /* execute1.vhdl:1103:29  */
  assign n11562_o = n9139_o[341];
  /* execute1.vhdl:1103:38  */
  assign n11563_o = ~n11562_o;
  /* execute1.vhdl:1104:59  */
  assign n11564_o = c_in[63:61];
  /* execute1.vhdl:1105:59  */
  assign n11565_o = c_in[59:32];
  assign n11566_o = ctrl[187:160];
  /* execute1.vhdl:1103:21  */
  assign n11567_o = n11563_o ? n11565_o : n11566_o;
  assign n11568_o = ctrl[191:189];
  /* execute1.vhdl:1103:21  */
  assign n11569_o = n11563_o ? n11564_o : n11568_o;
  /* execute1.vhdl:1109:28  */
  assign n11572_o = c_in[14];
  assign n11576_o = {1'b1, 1'b1};
  assign n11577_o = c_in[5:4];
  /* execute1.vhdl:1109:21  */
  assign n11578_o = n11572_o ? n11576_o : n11577_o;
  assign n11579_o = c_in[15];
  /* execute1.vhdl:1109:21  */
  assign n11580_o = n11572_o ? 1'b1 : n11579_o;
  assign n11581_o = c_in[11:6];
  assign n11582_o = c_in[3:1];
  assign n11583_o = c_in[31:16];
  assign n11584_o = c_in[14:13];
  /* execute1.vhdl:1115:54  */
  assign n11585_o = n9141_o[1];
  /* execute1.vhdl:1116:53  */
  assign n11586_o = c_in[11];
  /* execute1.vhdl:1116:70  */
  assign n11587_o = c_in[8];
  /* execute1.vhdl:1116:63  */
  assign n11588_o = n11586_o | n11587_o;
  /* execute1.vhdl:1115:64  */
  assign n11589_o = n11585_o & n11588_o;
  assign n11590_o = {n11581_o, n11578_o, n11582_o};
  assign n11591_o = {n11567_o, n11583_o, n11580_o, n11584_o};
  assign n11592_o = n11590_o[0];
  /* execute1.vhdl:1096:17  */
  assign n11593_o = n11559_o ? n11561_o : n11592_o;
  assign n11594_o = n11590_o[10:1];
  assign n11595_o = ctrl[139:130];
  /* execute1.vhdl:1096:17  */
  assign n11596_o = n11559_o ? n11595_o : n11594_o;
  assign n11597_o = n11591_o[1:0];
  assign n11598_o = ctrl[142:141];
  /* execute1.vhdl:1096:17  */
  assign n11599_o = n11559_o ? n11598_o : n11597_o;
  assign n11600_o = n11591_o[2];
  /* execute1.vhdl:1096:17  */
  assign n11601_o = n11559_o ? n11560_o : n11600_o;
  assign n11602_o = n11591_o[46:3];
  assign n11603_o = ctrl[187:144];
  /* execute1.vhdl:1096:17  */
  assign n11604_o = n11559_o ? n11603_o : n11602_o;
  assign n11605_o = ctrl[191:189];
  /* execute1.vhdl:1096:17  */
  assign n11606_o = n11559_o ? n11605_o : n11569_o;
  assign n11607_o = r[749];
  /* execute1.vhdl:1096:17  */
  assign n11608_o = n11559_o ? n11607_o : n11589_o;
  /* execute1.vhdl:1095:13  */
  assign n11610_o = n11096_o == 6'b100111;
  /* execute1.vhdl:1122:37  */
  assign n11612_o = n9139_o[83:77];
  /* common.vhdl:775:17  */
  assign n11617_o = n11612_o[5];
  /* execute1.vhdl:1123:44  */
  assign n11619_o = n9139_o[374:343];
  /* common.vhdl:708:40  */
  assign n11624_o = n11619_o[15:11];
  /* common.vhdl:708:61  */
  assign n11625_o = n11619_o[20:16];
  /* common.vhdl:708:55  */
  assign n11626_o = {n11624_o, n11625_o};
  /* execute1.vhdl:1123:50  */
  assign n11628_o = {22'b0, n11626_o};  //  uext
  /* execute1.vhdl:1123:50  */
  assign n11630_o = n11628_o == 32'b00000000000000000000000000000001;
  /* execute1.vhdl:1124:44  */
  assign n11631_o = c_in[31];
  /* execute1.vhdl:1125:44  */
  assign n11632_o = c_in[30];
  /* execute1.vhdl:1126:44  */
  assign n11633_o = c_in[29];
  /* execute1.vhdl:1127:46  */
  assign n11634_o = c_in[19];
  /* execute1.vhdl:1128:46  */
  assign n11635_o = c_in[18];
  assign n11636_o = {n11631_o, n11634_o, n11632_o, n11635_o, n11633_o};
  /* execute1.vhdl:1122:17  */
  assign n11637_o = n11731_o ? n11636_o : xerc_in;
  /* execute1.vhdl:1132:46  */
  assign n11639_o = n9139_o[374:343];
  /* common.vhdl:708:40  */
  assign n11644_o = n11639_o[15:11];
  /* common.vhdl:708:61  */
  assign n11645_o = n11639_o[20:16];
  /* common.vhdl:708:55  */
  assign n11646_o = {n11644_o, n11645_o};
  /* execute1.vhdl:1133:21  */
  assign n11649_o = n11646_o == 10'b0000010110;
  /* execute1.vhdl:1136:47  */
  assign n11650_o = c_in[31:0];
  /* execute1.vhdl:1135:21  */
  assign n11652_o = n11646_o == 10'b1011010100;
  /* execute1.vhdl:1137:21  */
  assign n11655_o = n11646_o == 10'b1100000011;
  /* execute1.vhdl:1137:36  */
  assign n11657_o = n11646_o == 10'b1100000100;
  /* execute1.vhdl:1137:36  */
  assign n11658_o = n11655_o | n11657_o;
  /* execute1.vhdl:1137:48  */
  assign n11660_o = n11646_o == 10'b1100000101;
  /* execute1.vhdl:1137:48  */
  assign n11661_o = n11658_o | n11660_o;
  /* execute1.vhdl:1137:60  */
  assign n11663_o = n11646_o == 10'b1100000110;
  /* execute1.vhdl:1137:60  */
  assign n11664_o = n11661_o | n11663_o;
  /* execute1.vhdl:1137:72  */
  assign n11666_o = n11646_o == 10'b1100000111;
  /* execute1.vhdl:1137:72  */
  assign n11667_o = n11664_o | n11666_o;
  /* execute1.vhdl:1137:84  */
  assign n11669_o = n11646_o == 10'b1100001000;
  /* execute1.vhdl:1137:84  */
  assign n11670_o = n11667_o | n11669_o;
  /* execute1.vhdl:1137:96  */
  assign n11672_o = n11646_o == 10'b1100001011;
  /* execute1.vhdl:1137:96  */
  assign n11673_o = n11670_o | n11672_o;
  /* execute1.vhdl:1138:36  */
  assign n11675_o = n11646_o == 10'b1100000001;
  /* execute1.vhdl:1138:36  */
  assign n11676_o = n11673_o | n11675_o;
  /* execute1.vhdl:1138:49  */
  assign n11678_o = n11646_o == 10'b1100000010;
  /* execute1.vhdl:1138:49  */
  assign n11679_o = n11676_o | n11678_o;
  /* execute1.vhdl:1138:62  */
  assign n11681_o = n11646_o == 10'b1100010011;
  /* execute1.vhdl:1138:62  */
  assign n11682_o = n11679_o | n11681_o;
  /* execute1.vhdl:1139:34  */
  assign n11684_o = n11646_o == 10'b1100010100;
  /* execute1.vhdl:1139:34  */
  assign n11685_o = n11682_o | n11684_o;
  /* execute1.vhdl:1139:45  */
  assign n11687_o = n11646_o == 10'b1100010101;
  /* execute1.vhdl:1139:45  */
  assign n11688_o = n11685_o | n11687_o;
  /* execute1.vhdl:1139:56  */
  assign n11690_o = n11646_o == 10'b1100010110;
  /* execute1.vhdl:1139:56  */
  assign n11691_o = n11688_o | n11690_o;
  /* execute1.vhdl:1139:67  */
  assign n11693_o = n11646_o == 10'b1100010111;
  /* execute1.vhdl:1139:67  */
  assign n11694_o = n11691_o | n11693_o;
  /* execute1.vhdl:1139:78  */
  assign n11696_o = n11646_o == 10'b1100011000;
  /* execute1.vhdl:1139:78  */
  assign n11697_o = n11694_o | n11696_o;
  /* execute1.vhdl:1139:89  */
  assign n11699_o = n11646_o == 10'b1100011011;
  /* execute1.vhdl:1139:89  */
  assign n11700_o = n11697_o | n11699_o;
  /* execute1.vhdl:1140:35  */
  assign n11702_o = n11646_o == 10'b1100011110;
  /* execute1.vhdl:1140:35  */
  assign n11703_o = n11700_o | n11702_o;
  /* execute1.vhdl:1140:47  */
  assign n11705_o = n11646_o == 10'b1100010001;
  /* execute1.vhdl:1140:47  */
  assign n11706_o = n11703_o | n11705_o;
  /* execute1.vhdl:1140:59  */
  assign n11708_o = n11646_o == 10'b1100010010;
  /* execute1.vhdl:1140:59  */
  assign n11709_o = n11706_o | n11708_o;
  /* execute1.vhdl:1140:71  */
  assign n11711_o = n11646_o == 10'b1100010000;
  /* execute1.vhdl:1140:71  */
  assign n11712_o = n11709_o | n11711_o;
  /* execute1.vhdl:1140:82  */
  assign n11714_o = n11646_o == 10'b1100011100;
  /* execute1.vhdl:1140:82  */
  assign n11715_o = n11712_o | n11714_o;
  /* execute1.vhdl:1140:93  */
  assign n11717_o = n11646_o == 10'b1100011101;
  /* execute1.vhdl:1140:93  */
  assign n11718_o = n11715_o | n11717_o;
  /* execute1.vhdl:1145:36  */
  assign n11719_o = ctrl[142];
  /* execute1.vhdl:1145:25  */
  assign n11722_o = n11719_o ? 1'b1 : 1'b0;
  assign n11723_o = {n11718_o, n11652_o, n11649_o};
  /* execute1.vhdl:1132:21  */
  always @*
    case (n11723_o)
      3'b100: n11724_o = n10752_o;
      3'b010: n11724_o = n10752_o;
      3'b001: n11724_o = c_in;
      default: n11724_o = n10752_o;
    endcase
  /* execute1.vhdl:1132:21  */
  always @*
    case (n11723_o)
      3'b100: n11725_o = 1'b1;
      3'b010: n11725_o = 1'b0;
      3'b001: n11725_o = 1'b0;
      default: n11725_o = 1'b0;
    endcase
  /* execute1.vhdl:1132:21  */
  always @*
    case (n11723_o)
      3'b100: n11726_o = n10737_o;
      3'b010: n11726_o = n11650_o;
      3'b001: n11726_o = n10737_o;
      default: n11726_o = n10737_o;
    endcase
  /* execute1.vhdl:1132:21  */
  always @*
    case (n11723_o)
      3'b100: n11728_o = 1'b0;
      3'b010: n11728_o = 1'b0;
      3'b001: n11728_o = 1'b0;
      default: n11728_o = n11722_o;
    endcase
  /* execute1.vhdl:1122:17  */
  assign n11729_o = n11617_o ? n10752_o : n11724_o;
  /* execute1.vhdl:1122:17  */
  assign n11730_o = n11617_o ? 1'b0 : n11725_o;
  /* execute1.vhdl:1122:17  */
  assign n11731_o = n11617_o & n11630_o;
  /* execute1.vhdl:1122:17  */
  assign n11732_o = n11617_o ? n10737_o : n11726_o;
  /* execute1.vhdl:1122:17  */
  assign n11734_o = n11617_o ? 1'b0 : n11728_o;
  /* execute1.vhdl:1119:13  */
  assign n11736_o = n11096_o == 6'b101000;
  /* execute1.vhdl:1151:25  */
  assign n11737_o = n9139_o[337];
  assign n11739_o = {n10737_o, 1'b0, 1'b0, n11032_o, n11086_o, n11081_o, 1'b0, 1'b0, 1'b0, 1'b0, n10837_o, n10836_o, n11068_o, n11071_o, 1'b0, n11065_o, n10834_o, n10817_o, n11056_o, n11031_o, n11059_o, n11027_o, n11053_o, n11023_o, n11047_o, n11019_o, n11041_o, n11015_o, n10823_o, n10822_o, n10715_o, n10815_o, n11011_o, n10816_o, xerc_in, n10826_o, n10825_o, n10829_o, n10828_o, 1'b1};
  assign n11743_o = n11739_o[119:0];
  assign n11744_o = n11739_o[353:122];
  assign n11745_o = {n11744_o, rotator_carry, rotator_carry, n11743_o};
  assign n11746_o = {n10817_o, n11056_o, n11031_o, n11059_o, n11027_o, n11053_o, n11023_o, n11047_o, n11019_o, n11041_o, n11015_o, n10823_o, n10822_o, n10715_o, n10815_o, n11011_o, n10816_o, xerc_in, n10826_o, n10825_o, n10829_o, n10828_o, 1'b1};
  /* execute1.vhdl:1151:17  */
  assign n11747_o = n11737_o ? n11745_o : n11746_o;
  /* execute1.vhdl:1150:13  */
  assign n11749_o = n11096_o == 6'b110000;
  /* execute1.vhdl:1150:25  */
  assign n11751_o = n11096_o == 6'b110001;
  /* execute1.vhdl:1150:25  */
  assign n11752_o = n11749_o | n11751_o;
  /* execute1.vhdl:1150:35  */
  assign n11754_o = n11096_o == 6'b110010;
  /* execute1.vhdl:1150:35  */
  assign n11755_o = n11752_o | n11754_o;
  /* execute1.vhdl:1150:45  */
  assign n11757_o = n11096_o == 6'b110101;
  /* execute1.vhdl:1150:45  */
  assign n11758_o = n11755_o | n11757_o;
  /* execute1.vhdl:1150:54  */
  assign n11760_o = n11096_o == 6'b110110;
  /* execute1.vhdl:1150:54  */
  assign n11761_o = n11758_o | n11760_o;
  /* execute1.vhdl:1150:63  */
  assign n11763_o = n11096_o == 6'b011000;
  /* execute1.vhdl:1150:63  */
  assign n11764_o = n11761_o | n11763_o;
  /* execute1.vhdl:1154:13  */
  assign n11766_o = n11096_o == 6'b110100;
  /* execute1.vhdl:1156:13  */
  assign n11770_o = n11096_o == 6'b011110;
  /* execute1.vhdl:1160:13  */
  assign n11772_o = n11096_o == 6'b011011;
  /* execute1.vhdl:1163:13  */
  assign n11778_o = n11096_o == 6'b101001;
  /* execute1.vhdl:1163:29  */
  assign n11780_o = n11096_o == 6'b101010;
  /* execute1.vhdl:1163:29  */
  assign n11781_o = n11778_o | n11780_o;
  /* execute1.vhdl:1163:42  */
  assign n11783_o = n11096_o == 6'b101011;
  /* execute1.vhdl:1163:42  */
  assign n11784_o = n11781_o | n11783_o;
  /* execute1.vhdl:1179:13  */
  assign n11790_o = n11096_o == 6'b010101;
  /* execute1.vhdl:1179:25  */
  assign n11792_o = n11096_o == 6'b010110;
  /* execute1.vhdl:1179:25  */
  assign n11793_o = n11790_o | n11792_o;
  /* execute1.vhdl:1179:35  */
  assign n11795_o = n11096_o == 6'b100101;
  /* execute1.vhdl:1179:35  */
  assign n11796_o = n11793_o | n11795_o;
  assign n11798_o = {n11796_o, n11784_o, n11772_o, n11770_o, n11766_o, n11764_o, n11736_o, n11610_o, n11558_o, n11556_o, n11554_o, n11364_o, n11362_o, n11360_o, n11358_o, n11356_o, n11354_o, n11346_o, n11312_o, n11230_o, n11223_o, n11200_o, n11198_o, n11196_o, n11194_o, n11179_o, n11177_o, n11136_o, n11119_o, n11109_o, n11098_o};
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11801_o = 1'b0;
      31'b0100000000000000000000000000000: n11801_o = 1'b0;
      31'b0010000000000000000000000000000: n11801_o = 1'b1;
      31'b0001000000000000000000000000000: n11801_o = 1'b0;
      31'b0000100000000000000000000000000: n11801_o = 1'b0;
      31'b0000010000000000000000000000000: n11801_o = 1'b0;
      31'b0000001000000000000000000000000: n11801_o = 1'b0;
      31'b0000000100000000000000000000000: n11801_o = 1'b0;
      31'b0000000010000000000000000000000: n11801_o = 1'b0;
      31'b0000000001000000000000000000000: n11801_o = 1'b0;
      31'b0000000000100000000000000000000: n11801_o = 1'b0;
      31'b0000000000010000000000000000000: n11801_o = 1'b0;
      31'b0000000000001000000000000000000: n11801_o = 1'b0;
      31'b0000000000000100000000000000000: n11801_o = 1'b0;
      31'b0000000000000010000000000000000: n11801_o = 1'b0;
      31'b0000000000000001000000000000000: n11801_o = 1'b0;
      31'b0000000000000000100000000000000: n11801_o = 1'b0;
      31'b0000000000000000010000000000000: n11801_o = 1'b0;
      31'b0000000000000000001000000000000: n11801_o = 1'b0;
      31'b0000000000000000000100000000000: n11801_o = 1'b0;
      31'b0000000000000000000010000000000: n11801_o = 1'b0;
      31'b0000000000000000000001000000000: n11801_o = 1'b0;
      31'b0000000000000000000000100000000: n11801_o = 1'b0;
      31'b0000000000000000000000010000000: n11801_o = 1'b0;
      31'b0000000000000000000000001000000: n11801_o = 1'b0;
      31'b0000000000000000000000000100000: n11801_o = 1'b0;
      31'b0000000000000000000000000010000: n11801_o = 1'b0;
      31'b0000000000000000000000000001000: n11801_o = 1'b0;
      31'b0000000000000000000000000000100: n11801_o = 1'b0;
      31'b0000000000000000000000000000010: n11801_o = 1'b0;
      31'b0000000000000000000000000000001: n11801_o = 1'b0;
      default: n11801_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11802_o = n10752_o;
      31'b0100000000000000000000000000000: n11802_o = n10752_o;
      31'b0010000000000000000000000000000: n11802_o = n10752_o;
      31'b0001000000000000000000000000000: n11802_o = n10752_o;
      31'b0000100000000000000000000000000: n11802_o = n10752_o;
      31'b0000010000000000000000000000000: n11802_o = n10752_o;
      31'b0000001000000000000000000000000: n11802_o = n11729_o;
      31'b0000000100000000000000000000000: n11802_o = n10752_o;
      31'b0000000010000000000000000000000: n11802_o = n10752_o;
      31'b0000000001000000000000000000000: n11802_o = n10752_o;
      31'b0000000000100000000000000000000: n11802_o = n10752_o;
      31'b0000000000010000000000000000000: n11802_o = n10752_o;
      31'b0000000000001000000000000000000: n11802_o = n10752_o;
      31'b0000000000000100000000000000000: n11802_o = n10752_o;
      31'b0000000000000010000000000000000: n11802_o = n10752_o;
      31'b0000000000000001000000000000000: n11802_o = n10752_o;
      31'b0000000000000000100000000000000: n11802_o = n10752_o;
      31'b0000000000000000010000000000000: n11802_o = n10752_o;
      31'b0000000000000000001000000000000: n11802_o = n10752_o;
      31'b0000000000000000000100000000000: n11802_o = n10752_o;
      31'b0000000000000000000010000000000: n11802_o = n10752_o;
      31'b0000000000000000000001000000000: n11802_o = n10752_o;
      31'b0000000000000000000000100000000: n11802_o = n10752_o;
      31'b0000000000000000000000010000000: n11802_o = n10752_o;
      31'b0000000000000000000000001000000: n11802_o = n10752_o;
      31'b0000000000000000000000000100000: n11802_o = n10752_o;
      31'b0000000000000000000000000010000: n11802_o = n10752_o;
      31'b0000000000000000000000000001000: n11802_o = n10752_o;
      31'b0000000000000000000000000000100: n11802_o = n10752_o;
      31'b0000000000000000000000000000010: n11802_o = n10752_o;
      31'b0000000000000000000000000000001: n11802_o = n10752_o;
      default: n11802_o = n10752_o;
    endcase
  assign n11803_o = n11338_o[0];
  assign n11804_o = ctrl[128];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11805_o = n11804_o;
      31'b0100000000000000000000000000000: n11805_o = n11804_o;
      31'b0010000000000000000000000000000: n11805_o = n11804_o;
      31'b0001000000000000000000000000000: n11805_o = n11804_o;
      31'b0000100000000000000000000000000: n11805_o = n11804_o;
      31'b0000010000000000000000000000000: n11805_o = n11804_o;
      31'b0000001000000000000000000000000: n11805_o = n11804_o;
      31'b0000000100000000000000000000000: n11805_o = n11804_o;
      31'b0000000010000000000000000000000: n11805_o = n11804_o;
      31'b0000000001000000000000000000000: n11805_o = n11804_o;
      31'b0000000000100000000000000000000: n11805_o = n11804_o;
      31'b0000000000010000000000000000000: n11805_o = n11804_o;
      31'b0000000000001000000000000000000: n11805_o = n11804_o;
      31'b0000000000000100000000000000000: n11805_o = n11804_o;
      31'b0000000000000010000000000000000: n11805_o = n11804_o;
      31'b0000000000000001000000000000000: n11805_o = n11804_o;
      31'b0000000000000000100000000000000: n11805_o = n11804_o;
      31'b0000000000000000010000000000000: n11805_o = n11803_o;
      31'b0000000000000000001000000000000: n11805_o = n11804_o;
      31'b0000000000000000000100000000000: n11805_o = n11804_o;
      31'b0000000000000000000010000000000: n11805_o = n11804_o;
      31'b0000000000000000000001000000000: n11805_o = n11804_o;
      31'b0000000000000000000000100000000: n11805_o = n11804_o;
      31'b0000000000000000000000010000000: n11805_o = n11804_o;
      31'b0000000000000000000000001000000: n11805_o = n11804_o;
      31'b0000000000000000000000000100000: n11805_o = n11804_o;
      31'b0000000000000000000000000010000: n11805_o = n11804_o;
      31'b0000000000000000000000000001000: n11805_o = n11804_o;
      31'b0000000000000000000000000000100: n11805_o = n11804_o;
      31'b0000000000000000000000000000010: n11805_o = n11804_o;
      31'b0000000000000000000000000000001: n11805_o = n11804_o;
      default: n11805_o = n11804_o;
    endcase
  assign n11806_o = n11338_o[1];
  assign n11807_o = ctrl[129];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11808_o = n11807_o;
      31'b0100000000000000000000000000000: n11808_o = n11807_o;
      31'b0010000000000000000000000000000: n11808_o = n11807_o;
      31'b0001000000000000000000000000000: n11808_o = n11807_o;
      31'b0000100000000000000000000000000: n11808_o = n11807_o;
      31'b0000010000000000000000000000000: n11808_o = n11807_o;
      31'b0000001000000000000000000000000: n11808_o = n11807_o;
      31'b0000000100000000000000000000000: n11808_o = n11593_o;
      31'b0000000010000000000000000000000: n11808_o = n11807_o;
      31'b0000000001000000000000000000000: n11808_o = n11807_o;
      31'b0000000000100000000000000000000: n11808_o = n11807_o;
      31'b0000000000010000000000000000000: n11808_o = n11807_o;
      31'b0000000000001000000000000000000: n11808_o = n11807_o;
      31'b0000000000000100000000000000000: n11808_o = n11807_o;
      31'b0000000000000010000000000000000: n11808_o = n11807_o;
      31'b0000000000000001000000000000000: n11808_o = n11807_o;
      31'b0000000000000000100000000000000: n11808_o = n11807_o;
      31'b0000000000000000010000000000000: n11808_o = n11806_o;
      31'b0000000000000000001000000000000: n11808_o = n11807_o;
      31'b0000000000000000000100000000000: n11808_o = n11807_o;
      31'b0000000000000000000010000000000: n11808_o = n11807_o;
      31'b0000000000000000000001000000000: n11808_o = n11807_o;
      31'b0000000000000000000000100000000: n11808_o = n11807_o;
      31'b0000000000000000000000010000000: n11808_o = n11807_o;
      31'b0000000000000000000000001000000: n11808_o = n11807_o;
      31'b0000000000000000000000000100000: n11808_o = n11807_o;
      31'b0000000000000000000000000010000: n11808_o = n11807_o;
      31'b0000000000000000000000000001000: n11808_o = n11807_o;
      31'b0000000000000000000000000000100: n11808_o = n11807_o;
      31'b0000000000000000000000000000010: n11808_o = n11807_o;
      31'b0000000000000000000000000000001: n11808_o = n11807_o;
      default: n11808_o = n11807_o;
    endcase
  assign n11809_o = n11338_o[3:2];
  assign n11810_o = n11596_o[1:0];
  assign n11811_o = ctrl[131:130];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11812_o = n11811_o;
      31'b0100000000000000000000000000000: n11812_o = n11811_o;
      31'b0010000000000000000000000000000: n11812_o = n11811_o;
      31'b0001000000000000000000000000000: n11812_o = n11811_o;
      31'b0000100000000000000000000000000: n11812_o = n11811_o;
      31'b0000010000000000000000000000000: n11812_o = n11811_o;
      31'b0000001000000000000000000000000: n11812_o = n11811_o;
      31'b0000000100000000000000000000000: n11812_o = n11810_o;
      31'b0000000010000000000000000000000: n11812_o = n11811_o;
      31'b0000000001000000000000000000000: n11812_o = n11811_o;
      31'b0000000000100000000000000000000: n11812_o = n11811_o;
      31'b0000000000010000000000000000000: n11812_o = n11811_o;
      31'b0000000000001000000000000000000: n11812_o = n11811_o;
      31'b0000000000000100000000000000000: n11812_o = n11811_o;
      31'b0000000000000010000000000000000: n11812_o = n11811_o;
      31'b0000000000000001000000000000000: n11812_o = n11811_o;
      31'b0000000000000000100000000000000: n11812_o = n11811_o;
      31'b0000000000000000010000000000000: n11812_o = n11809_o;
      31'b0000000000000000001000000000000: n11812_o = n11811_o;
      31'b0000000000000000000100000000000: n11812_o = n11811_o;
      31'b0000000000000000000010000000000: n11812_o = n11811_o;
      31'b0000000000000000000001000000000: n11812_o = n11811_o;
      31'b0000000000000000000000100000000: n11812_o = n11811_o;
      31'b0000000000000000000000010000000: n11812_o = n11811_o;
      31'b0000000000000000000000001000000: n11812_o = n11811_o;
      31'b0000000000000000000000000100000: n11812_o = n11811_o;
      31'b0000000000000000000000000010000: n11812_o = n11811_o;
      31'b0000000000000000000000000001000: n11812_o = n11811_o;
      31'b0000000000000000000000000000100: n11812_o = n11811_o;
      31'b0000000000000000000000000000010: n11812_o = n11811_o;
      31'b0000000000000000000000000000001: n11812_o = n11811_o;
      default: n11812_o = n11811_o;
    endcase
  assign n11813_o = n11596_o[3:2];
  assign n11814_o = ctrl[133:132];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11815_o = n11814_o;
      31'b0100000000000000000000000000000: n11815_o = n11814_o;
      31'b0010000000000000000000000000000: n11815_o = n11814_o;
      31'b0001000000000000000000000000000: n11815_o = n11814_o;
      31'b0000100000000000000000000000000: n11815_o = n11814_o;
      31'b0000010000000000000000000000000: n11815_o = n11814_o;
      31'b0000001000000000000000000000000: n11815_o = n11814_o;
      31'b0000000100000000000000000000000: n11815_o = n11813_o;
      31'b0000000010000000000000000000000: n11815_o = n11814_o;
      31'b0000000001000000000000000000000: n11815_o = n11814_o;
      31'b0000000000100000000000000000000: n11815_o = n11814_o;
      31'b0000000000010000000000000000000: n11815_o = n11814_o;
      31'b0000000000001000000000000000000: n11815_o = n11814_o;
      31'b0000000000000100000000000000000: n11815_o = n11814_o;
      31'b0000000000000010000000000000000: n11815_o = n11814_o;
      31'b0000000000000001000000000000000: n11815_o = n11814_o;
      31'b0000000000000000100000000000000: n11815_o = n11814_o;
      31'b0000000000000000010000000000000: n11815_o = n11334_o;
      31'b0000000000000000001000000000000: n11815_o = n11814_o;
      31'b0000000000000000000100000000000: n11815_o = n11814_o;
      31'b0000000000000000000010000000000: n11815_o = n11814_o;
      31'b0000000000000000000001000000000: n11815_o = n11814_o;
      31'b0000000000000000000000100000000: n11815_o = n11814_o;
      31'b0000000000000000000000010000000: n11815_o = n11814_o;
      31'b0000000000000000000000001000000: n11815_o = n11814_o;
      31'b0000000000000000000000000100000: n11815_o = n11814_o;
      31'b0000000000000000000000000010000: n11815_o = n11814_o;
      31'b0000000000000000000000000001000: n11815_o = n11814_o;
      31'b0000000000000000000000000000100: n11815_o = n11814_o;
      31'b0000000000000000000000000000010: n11815_o = n11814_o;
      31'b0000000000000000000000000000001: n11815_o = n11814_o;
      default: n11815_o = n11814_o;
    endcase
  assign n11816_o = n11339_o[5:0];
  assign n11817_o = n11596_o[9:4];
  assign n11818_o = ctrl[139:134];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11819_o = n11818_o;
      31'b0100000000000000000000000000000: n11819_o = n11818_o;
      31'b0010000000000000000000000000000: n11819_o = n11818_o;
      31'b0001000000000000000000000000000: n11819_o = n11818_o;
      31'b0000100000000000000000000000000: n11819_o = n11818_o;
      31'b0000010000000000000000000000000: n11819_o = n11818_o;
      31'b0000001000000000000000000000000: n11819_o = n11818_o;
      31'b0000000100000000000000000000000: n11819_o = n11817_o;
      31'b0000000010000000000000000000000: n11819_o = n11818_o;
      31'b0000000001000000000000000000000: n11819_o = n11818_o;
      31'b0000000000100000000000000000000: n11819_o = n11818_o;
      31'b0000000000010000000000000000000: n11819_o = n11818_o;
      31'b0000000000001000000000000000000: n11819_o = n11818_o;
      31'b0000000000000100000000000000000: n11819_o = n11818_o;
      31'b0000000000000010000000000000000: n11819_o = n11818_o;
      31'b0000000000000001000000000000000: n11819_o = n11818_o;
      31'b0000000000000000100000000000000: n11819_o = n11818_o;
      31'b0000000000000000010000000000000: n11819_o = n11816_o;
      31'b0000000000000000001000000000000: n11819_o = n11818_o;
      31'b0000000000000000000100000000000: n11819_o = n11818_o;
      31'b0000000000000000000010000000000: n11819_o = n11818_o;
      31'b0000000000000000000001000000000: n11819_o = n11818_o;
      31'b0000000000000000000000100000000: n11819_o = n11818_o;
      31'b0000000000000000000000010000000: n11819_o = n11818_o;
      31'b0000000000000000000000001000000: n11819_o = n11818_o;
      31'b0000000000000000000000000100000: n11819_o = n11818_o;
      31'b0000000000000000000000000010000: n11819_o = n11818_o;
      31'b0000000000000000000000000001000: n11819_o = n11818_o;
      31'b0000000000000000000000000000100: n11819_o = n11818_o;
      31'b0000000000000000000000000000010: n11819_o = n11818_o;
      31'b0000000000000000000000000000001: n11819_o = n11818_o;
      default: n11819_o = n11818_o;
    endcase
  assign n11820_o = n11339_o[6];
  assign n11821_o = ctrl[140];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11822_o = n11821_o;
      31'b0100000000000000000000000000000: n11822_o = n11821_o;
      31'b0010000000000000000000000000000: n11822_o = n11821_o;
      31'b0001000000000000000000000000000: n11822_o = n11821_o;
      31'b0000100000000000000000000000000: n11822_o = n11821_o;
      31'b0000010000000000000000000000000: n11822_o = n11821_o;
      31'b0000001000000000000000000000000: n11822_o = n11821_o;
      31'b0000000100000000000000000000000: n11822_o = n11821_o;
      31'b0000000010000000000000000000000: n11822_o = n11821_o;
      31'b0000000001000000000000000000000: n11822_o = n11821_o;
      31'b0000000000100000000000000000000: n11822_o = n11821_o;
      31'b0000000000010000000000000000000: n11822_o = n11821_o;
      31'b0000000000001000000000000000000: n11822_o = n11821_o;
      31'b0000000000000100000000000000000: n11822_o = n11821_o;
      31'b0000000000000010000000000000000: n11822_o = n11821_o;
      31'b0000000000000001000000000000000: n11822_o = n11821_o;
      31'b0000000000000000100000000000000: n11822_o = n11821_o;
      31'b0000000000000000010000000000000: n11822_o = n11820_o;
      31'b0000000000000000001000000000000: n11822_o = n11821_o;
      31'b0000000000000000000100000000000: n11822_o = n11821_o;
      31'b0000000000000000000010000000000: n11822_o = n11821_o;
      31'b0000000000000000000001000000000: n11822_o = n11821_o;
      31'b0000000000000000000000100000000: n11822_o = n11821_o;
      31'b0000000000000000000000010000000: n11822_o = n11821_o;
      31'b0000000000000000000000001000000: n11822_o = n11821_o;
      31'b0000000000000000000000000100000: n11822_o = n11821_o;
      31'b0000000000000000000000000010000: n11822_o = n11821_o;
      31'b0000000000000000000000000001000: n11822_o = n11821_o;
      31'b0000000000000000000000000000100: n11822_o = n11821_o;
      31'b0000000000000000000000000000010: n11822_o = n11821_o;
      31'b0000000000000000000000000000001: n11822_o = n11821_o;
      default: n11822_o = n11821_o;
    endcase
  assign n11823_o = n11339_o[8:7];
  assign n11824_o = ctrl[142:141];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11825_o = n11824_o;
      31'b0100000000000000000000000000000: n11825_o = n11824_o;
      31'b0010000000000000000000000000000: n11825_o = n11824_o;
      31'b0001000000000000000000000000000: n11825_o = n11824_o;
      31'b0000100000000000000000000000000: n11825_o = n11824_o;
      31'b0000010000000000000000000000000: n11825_o = n11824_o;
      31'b0000001000000000000000000000000: n11825_o = n11824_o;
      31'b0000000100000000000000000000000: n11825_o = n11599_o;
      31'b0000000010000000000000000000000: n11825_o = n11824_o;
      31'b0000000001000000000000000000000: n11825_o = n11824_o;
      31'b0000000000100000000000000000000: n11825_o = n11824_o;
      31'b0000000000010000000000000000000: n11825_o = n11824_o;
      31'b0000000000001000000000000000000: n11825_o = n11824_o;
      31'b0000000000000100000000000000000: n11825_o = n11824_o;
      31'b0000000000000010000000000000000: n11825_o = n11824_o;
      31'b0000000000000001000000000000000: n11825_o = n11824_o;
      31'b0000000000000000100000000000000: n11825_o = n11824_o;
      31'b0000000000000000010000000000000: n11825_o = n11823_o;
      31'b0000000000000000001000000000000: n11825_o = n11824_o;
      31'b0000000000000000000100000000000: n11825_o = n11824_o;
      31'b0000000000000000000010000000000: n11825_o = n11824_o;
      31'b0000000000000000000001000000000: n11825_o = n11824_o;
      31'b0000000000000000000000100000000: n11825_o = n11824_o;
      31'b0000000000000000000000010000000: n11825_o = n11824_o;
      31'b0000000000000000000000001000000: n11825_o = n11824_o;
      31'b0000000000000000000000000100000: n11825_o = n11824_o;
      31'b0000000000000000000000000010000: n11825_o = n11824_o;
      31'b0000000000000000000000000001000: n11825_o = n11824_o;
      31'b0000000000000000000000000000100: n11825_o = n11824_o;
      31'b0000000000000000000000000000010: n11825_o = n11824_o;
      31'b0000000000000000000000000000001: n11825_o = n11824_o;
      default: n11825_o = n11824_o;
    endcase
  assign n11826_o = ctrl[143];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11827_o = n11826_o;
      31'b0100000000000000000000000000000: n11827_o = n11826_o;
      31'b0010000000000000000000000000000: n11827_o = n11826_o;
      31'b0001000000000000000000000000000: n11827_o = n11826_o;
      31'b0000100000000000000000000000000: n11827_o = n11826_o;
      31'b0000010000000000000000000000000: n11827_o = n11826_o;
      31'b0000001000000000000000000000000: n11827_o = n11826_o;
      31'b0000000100000000000000000000000: n11827_o = n11601_o;
      31'b0000000010000000000000000000000: n11827_o = n11826_o;
      31'b0000000001000000000000000000000: n11827_o = n11826_o;
      31'b0000000000100000000000000000000: n11827_o = n11826_o;
      31'b0000000000010000000000000000000: n11827_o = n11826_o;
      31'b0000000000001000000000000000000: n11827_o = n11826_o;
      31'b0000000000000100000000000000000: n11827_o = n11826_o;
      31'b0000000000000010000000000000000: n11827_o = n11826_o;
      31'b0000000000000001000000000000000: n11827_o = n11826_o;
      31'b0000000000000000100000000000000: n11827_o = n11826_o;
      31'b0000000000000000010000000000000: n11827_o = n11336_o;
      31'b0000000000000000001000000000000: n11827_o = n11826_o;
      31'b0000000000000000000100000000000: n11827_o = n11826_o;
      31'b0000000000000000000010000000000: n11827_o = n11826_o;
      31'b0000000000000000000001000000000: n11827_o = n11826_o;
      31'b0000000000000000000000100000000: n11827_o = n11826_o;
      31'b0000000000000000000000010000000: n11827_o = n11826_o;
      31'b0000000000000000000000001000000: n11827_o = n11826_o;
      31'b0000000000000000000000000100000: n11827_o = n11826_o;
      31'b0000000000000000000000000010000: n11827_o = n11826_o;
      31'b0000000000000000000000000001000: n11827_o = n11826_o;
      31'b0000000000000000000000000000100: n11827_o = n11826_o;
      31'b0000000000000000000000000000010: n11827_o = n11826_o;
      31'b0000000000000000000000000000001: n11827_o = n11826_o;
      default: n11827_o = n11826_o;
    endcase
  assign n11828_o = n11604_o[5:0];
  assign n11829_o = ctrl[149:144];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11830_o = n11829_o;
      31'b0100000000000000000000000000000: n11830_o = n11829_o;
      31'b0010000000000000000000000000000: n11830_o = n11829_o;
      31'b0001000000000000000000000000000: n11830_o = n11829_o;
      31'b0000100000000000000000000000000: n11830_o = n11829_o;
      31'b0000010000000000000000000000000: n11830_o = n11829_o;
      31'b0000001000000000000000000000000: n11830_o = n11829_o;
      31'b0000000100000000000000000000000: n11830_o = n11828_o;
      31'b0000000010000000000000000000000: n11830_o = n11829_o;
      31'b0000000001000000000000000000000: n11830_o = n11829_o;
      31'b0000000000100000000000000000000: n11830_o = n11829_o;
      31'b0000000000010000000000000000000: n11830_o = n11829_o;
      31'b0000000000001000000000000000000: n11830_o = n11829_o;
      31'b0000000000000100000000000000000: n11830_o = n11829_o;
      31'b0000000000000010000000000000000: n11830_o = n11829_o;
      31'b0000000000000001000000000000000: n11830_o = n11829_o;
      31'b0000000000000000100000000000000: n11830_o = n11829_o;
      31'b0000000000000000010000000000000: n11830_o = n11829_o;
      31'b0000000000000000001000000000000: n11830_o = n11829_o;
      31'b0000000000000000000100000000000: n11830_o = n11829_o;
      31'b0000000000000000000010000000000: n11830_o = n11829_o;
      31'b0000000000000000000001000000000: n11830_o = n11829_o;
      31'b0000000000000000000000100000000: n11830_o = n11829_o;
      31'b0000000000000000000000010000000: n11830_o = n11829_o;
      31'b0000000000000000000000001000000: n11830_o = n11829_o;
      31'b0000000000000000000000000100000: n11830_o = n11829_o;
      31'b0000000000000000000000000010000: n11830_o = n11829_o;
      31'b0000000000000000000000000001000: n11830_o = n11829_o;
      31'b0000000000000000000000000000100: n11830_o = n11829_o;
      31'b0000000000000000000000000000010: n11830_o = n11829_o;
      31'b0000000000000000000000000000001: n11830_o = n11829_o;
      default: n11830_o = n11829_o;
    endcase
  assign n11831_o = n11604_o[10:6];
  assign n11832_o = ctrl[154:150];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11833_o = n11832_o;
      31'b0100000000000000000000000000000: n11833_o = n11832_o;
      31'b0010000000000000000000000000000: n11833_o = n11832_o;
      31'b0001000000000000000000000000000: n11833_o = n11832_o;
      31'b0000100000000000000000000000000: n11833_o = n11832_o;
      31'b0000010000000000000000000000000: n11833_o = n11832_o;
      31'b0000001000000000000000000000000: n11833_o = n11832_o;
      31'b0000000100000000000000000000000: n11833_o = n11831_o;
      31'b0000000010000000000000000000000: n11833_o = n11832_o;
      31'b0000000001000000000000000000000: n11833_o = n11832_o;
      31'b0000000000100000000000000000000: n11833_o = n11832_o;
      31'b0000000000010000000000000000000: n11833_o = n11832_o;
      31'b0000000000001000000000000000000: n11833_o = n11832_o;
      31'b0000000000000100000000000000000: n11833_o = n11832_o;
      31'b0000000000000010000000000000000: n11833_o = n11832_o;
      31'b0000000000000001000000000000000: n11833_o = n11832_o;
      31'b0000000000000000100000000000000: n11833_o = n11832_o;
      31'b0000000000000000010000000000000: n11833_o = n11326_o;
      31'b0000000000000000001000000000000: n11833_o = n11832_o;
      31'b0000000000000000000100000000000: n11833_o = n11832_o;
      31'b0000000000000000000010000000000: n11833_o = n11832_o;
      31'b0000000000000000000001000000000: n11833_o = n11832_o;
      31'b0000000000000000000000100000000: n11833_o = n11832_o;
      31'b0000000000000000000000010000000: n11833_o = n11832_o;
      31'b0000000000000000000000001000000: n11833_o = n11832_o;
      31'b0000000000000000000000000100000: n11833_o = n11832_o;
      31'b0000000000000000000000000010000: n11833_o = n11832_o;
      31'b0000000000000000000000000001000: n11833_o = n11832_o;
      31'b0000000000000000000000000000100: n11833_o = n11832_o;
      31'b0000000000000000000000000000010: n11833_o = n11832_o;
      31'b0000000000000000000000000000001: n11833_o = n11832_o;
      default: n11833_o = n11832_o;
    endcase
  assign n11834_o = n11604_o[14:11];
  assign n11835_o = ctrl[158:155];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11836_o = n11835_o;
      31'b0100000000000000000000000000000: n11836_o = n11835_o;
      31'b0010000000000000000000000000000: n11836_o = n11835_o;
      31'b0001000000000000000000000000000: n11836_o = n11835_o;
      31'b0000100000000000000000000000000: n11836_o = n11835_o;
      31'b0000010000000000000000000000000: n11836_o = n11835_o;
      31'b0000001000000000000000000000000: n11836_o = n11835_o;
      31'b0000000100000000000000000000000: n11836_o = n11834_o;
      31'b0000000010000000000000000000000: n11836_o = n11835_o;
      31'b0000000001000000000000000000000: n11836_o = n11835_o;
      31'b0000000000100000000000000000000: n11836_o = n11835_o;
      31'b0000000000010000000000000000000: n11836_o = n11835_o;
      31'b0000000000001000000000000000000: n11836_o = n11835_o;
      31'b0000000000000100000000000000000: n11836_o = n11835_o;
      31'b0000000000000010000000000000000: n11836_o = n11835_o;
      31'b0000000000000001000000000000000: n11836_o = n11835_o;
      31'b0000000000000000100000000000000: n11836_o = n11835_o;
      31'b0000000000000000010000000000000: n11836_o = n11835_o;
      31'b0000000000000000001000000000000: n11836_o = n11835_o;
      31'b0000000000000000000100000000000: n11836_o = n11835_o;
      31'b0000000000000000000010000000000: n11836_o = n11835_o;
      31'b0000000000000000000001000000000: n11836_o = n11835_o;
      31'b0000000000000000000000100000000: n11836_o = n11835_o;
      31'b0000000000000000000000010000000: n11836_o = n11835_o;
      31'b0000000000000000000000001000000: n11836_o = n11835_o;
      31'b0000000000000000000000000100000: n11836_o = n11835_o;
      31'b0000000000000000000000000010000: n11836_o = n11835_o;
      31'b0000000000000000000000000001000: n11836_o = n11835_o;
      31'b0000000000000000000000000000100: n11836_o = n11835_o;
      31'b0000000000000000000000000000010: n11836_o = n11835_o;
      31'b0000000000000000000000000000001: n11836_o = n11835_o;
      default: n11836_o = n11835_o;
    endcase
  assign n11837_o = n11325_o[28:0];
  assign n11838_o = n11604_o[43:15];
  assign n11839_o = ctrl[187:159];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11840_o = n11839_o;
      31'b0100000000000000000000000000000: n11840_o = n11839_o;
      31'b0010000000000000000000000000000: n11840_o = n11839_o;
      31'b0001000000000000000000000000000: n11840_o = n11839_o;
      31'b0000100000000000000000000000000: n11840_o = n11839_o;
      31'b0000010000000000000000000000000: n11840_o = n11839_o;
      31'b0000001000000000000000000000000: n11840_o = n11839_o;
      31'b0000000100000000000000000000000: n11840_o = n11838_o;
      31'b0000000010000000000000000000000: n11840_o = n11839_o;
      31'b0000000001000000000000000000000: n11840_o = n11839_o;
      31'b0000000000100000000000000000000: n11840_o = n11839_o;
      31'b0000000000010000000000000000000: n11840_o = n11839_o;
      31'b0000000000001000000000000000000: n11840_o = n11839_o;
      31'b0000000000000100000000000000000: n11840_o = n11839_o;
      31'b0000000000000010000000000000000: n11840_o = n11839_o;
      31'b0000000000000001000000000000000: n11840_o = n11839_o;
      31'b0000000000000000100000000000000: n11840_o = n11839_o;
      31'b0000000000000000010000000000000: n11840_o = n11837_o;
      31'b0000000000000000001000000000000: n11840_o = n11839_o;
      31'b0000000000000000000100000000000: n11840_o = n11839_o;
      31'b0000000000000000000010000000000: n11840_o = n11839_o;
      31'b0000000000000000000001000000000: n11840_o = n11839_o;
      31'b0000000000000000000000100000000: n11840_o = n11839_o;
      31'b0000000000000000000000010000000: n11840_o = n11839_o;
      31'b0000000000000000000000001000000: n11840_o = n11839_o;
      31'b0000000000000000000000000100000: n11840_o = n11839_o;
      31'b0000000000000000000000000010000: n11840_o = n11839_o;
      31'b0000000000000000000000000001000: n11840_o = n11839_o;
      31'b0000000000000000000000000000100: n11840_o = n11839_o;
      31'b0000000000000000000000000000010: n11840_o = n11839_o;
      31'b0000000000000000000000000000001: n11840_o = n11839_o;
      default: n11840_o = n11839_o;
    endcase
  assign n11841_o = n11325_o[29];
  assign n11842_o = ctrl[188];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11843_o = n11842_o;
      31'b0100000000000000000000000000000: n11843_o = n11842_o;
      31'b0010000000000000000000000000000: n11843_o = n11842_o;
      31'b0001000000000000000000000000000: n11843_o = n11842_o;
      31'b0000100000000000000000000000000: n11843_o = n11842_o;
      31'b0000010000000000000000000000000: n11843_o = n11842_o;
      31'b0000001000000000000000000000000: n11843_o = n11842_o;
      31'b0000000100000000000000000000000: n11843_o = n11842_o;
      31'b0000000010000000000000000000000: n11843_o = n11842_o;
      31'b0000000001000000000000000000000: n11843_o = n11842_o;
      31'b0000000000100000000000000000000: n11843_o = n11842_o;
      31'b0000000000010000000000000000000: n11843_o = n11842_o;
      31'b0000000000001000000000000000000: n11843_o = n11842_o;
      31'b0000000000000100000000000000000: n11843_o = n11842_o;
      31'b0000000000000010000000000000000: n11843_o = n11842_o;
      31'b0000000000000001000000000000000: n11843_o = n11842_o;
      31'b0000000000000000100000000000000: n11843_o = n11842_o;
      31'b0000000000000000010000000000000: n11843_o = n11841_o;
      31'b0000000000000000001000000000000: n11843_o = n11842_o;
      31'b0000000000000000000100000000000: n11843_o = n11842_o;
      31'b0000000000000000000010000000000: n11843_o = n11842_o;
      31'b0000000000000000000001000000000: n11843_o = n11842_o;
      31'b0000000000000000000000100000000: n11843_o = n11842_o;
      31'b0000000000000000000000010000000: n11843_o = n11842_o;
      31'b0000000000000000000000001000000: n11843_o = n11842_o;
      31'b0000000000000000000000000100000: n11843_o = n11842_o;
      31'b0000000000000000000000000010000: n11843_o = n11842_o;
      31'b0000000000000000000000000001000: n11843_o = n11842_o;
      31'b0000000000000000000000000000100: n11843_o = n11842_o;
      31'b0000000000000000000000000000010: n11843_o = n11842_o;
      31'b0000000000000000000000000000001: n11843_o = n11842_o;
      default: n11843_o = n11842_o;
    endcase
  assign n11844_o = n11325_o[32:30];
  assign n11845_o = ctrl[191:189];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11846_o = n11845_o;
      31'b0100000000000000000000000000000: n11846_o = n11845_o;
      31'b0010000000000000000000000000000: n11846_o = n11845_o;
      31'b0001000000000000000000000000000: n11846_o = n11845_o;
      31'b0000100000000000000000000000000: n11846_o = n11845_o;
      31'b0000010000000000000000000000000: n11846_o = n11845_o;
      31'b0000001000000000000000000000000: n11846_o = n11845_o;
      31'b0000000100000000000000000000000: n11846_o = n11606_o;
      31'b0000000010000000000000000000000: n11846_o = n11845_o;
      31'b0000000001000000000000000000000: n11846_o = n11845_o;
      31'b0000000000100000000000000000000: n11846_o = n11845_o;
      31'b0000000000010000000000000000000: n11846_o = n11845_o;
      31'b0000000000001000000000000000000: n11846_o = n11845_o;
      31'b0000000000000100000000000000000: n11846_o = n11845_o;
      31'b0000000000000010000000000000000: n11846_o = n11845_o;
      31'b0000000000000001000000000000000: n11846_o = n11845_o;
      31'b0000000000000000100000000000000: n11846_o = n11845_o;
      31'b0000000000000000010000000000000: n11846_o = n11844_o;
      31'b0000000000000000001000000000000: n11846_o = n11845_o;
      31'b0000000000000000000100000000000: n11846_o = n11845_o;
      31'b0000000000000000000010000000000: n11846_o = n11845_o;
      31'b0000000000000000000001000000000: n11846_o = n11845_o;
      31'b0000000000000000000000100000000: n11846_o = n11845_o;
      31'b0000000000000000000000010000000: n11846_o = n11845_o;
      31'b0000000000000000000000001000000: n11846_o = n11845_o;
      31'b0000000000000000000000000100000: n11846_o = n11845_o;
      31'b0000000000000000000000000010000: n11846_o = n11845_o;
      31'b0000000000000000000000000001000: n11846_o = n11845_o;
      31'b0000000000000000000000000000100: n11846_o = n11845_o;
      31'b0000000000000000000000000000010: n11846_o = n11845_o;
      31'b0000000000000000000000000000001: n11846_o = n11845_o;
      default: n11846_o = n11845_o;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0100000000000000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0010000000000000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0001000000000000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000100000000000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000010000000000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000001000000000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000100000000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000010000000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000001000000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000100000000000000000000: n11848_o = n11552_o;
      31'b0000000000010000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000001000000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000100000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000010000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000001000000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000100000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000010000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000001000000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000100000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000010000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000001000000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000000100000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000000010000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000000001000000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000000000100000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000000000010000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000000000001000: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000000000000100: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000000000000010: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      31'b0000000000000000000000000000001: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
      default: n11848_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11849_o = 1'b0;
      31'b0100000000000000000000000000000: n11849_o = 1'b1;
      31'b0010000000000000000000000000000: n11849_o = 1'b0;
      31'b0001000000000000000000000000000: n11849_o = 1'b0;
      31'b0000100000000000000000000000000: n11849_o = 1'b0;
      31'b0000010000000000000000000000000: n11849_o = 1'b0;
      31'b0000001000000000000000000000000: n11849_o = 1'b0;
      31'b0000000100000000000000000000000: n11849_o = 1'b0;
      31'b0000000010000000000000000000000: n11849_o = 1'b0;
      31'b0000000001000000000000000000000: n11849_o = 1'b0;
      31'b0000000000100000000000000000000: n11849_o = 1'b0;
      31'b0000000000010000000000000000000: n11849_o = 1'b0;
      31'b0000000000001000000000000000000: n11849_o = 1'b0;
      31'b0000000000000100000000000000000: n11849_o = 1'b0;
      31'b0000000000000010000000000000000: n11849_o = 1'b0;
      31'b0000000000000001000000000000000: n11849_o = 1'b0;
      31'b0000000000000000100000000000000: n11849_o = 1'b0;
      31'b0000000000000000010000000000000: n11849_o = 1'b0;
      31'b0000000000000000001000000000000: n11849_o = 1'b0;
      31'b0000000000000000000100000000000: n11849_o = 1'b0;
      31'b0000000000000000000010000000000: n11849_o = 1'b0;
      31'b0000000000000000000001000000000: n11849_o = 1'b0;
      31'b0000000000000000000000100000000: n11849_o = 1'b0;
      31'b0000000000000000000000010000000: n11849_o = 1'b0;
      31'b0000000000000000000000001000000: n11849_o = 1'b0;
      31'b0000000000000000000000000100000: n11849_o = 1'b0;
      31'b0000000000000000000000000010000: n11849_o = 1'b0;
      31'b0000000000000000000000000001000: n11849_o = 1'b0;
      31'b0000000000000000000000000000100: n11849_o = 1'b0;
      31'b0000000000000000000000000000010: n11849_o = 1'b0;
      31'b0000000000000000000000000000001: n11849_o = 1'b0;
      default: n11849_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11850_o = 1'b1;
      31'b0100000000000000000000000000000: n11850_o = 1'b0;
      31'b0010000000000000000000000000000: n11850_o = 1'b0;
      31'b0001000000000000000000000000000: n11850_o = 1'b0;
      31'b0000100000000000000000000000000: n11850_o = 1'b0;
      31'b0000010000000000000000000000000: n11850_o = 1'b0;
      31'b0000001000000000000000000000000: n11850_o = 1'b0;
      31'b0000000100000000000000000000000: n11850_o = 1'b0;
      31'b0000000010000000000000000000000: n11850_o = 1'b0;
      31'b0000000001000000000000000000000: n11850_o = 1'b0;
      31'b0000000000100000000000000000000: n11850_o = 1'b0;
      31'b0000000000010000000000000000000: n11850_o = 1'b0;
      31'b0000000000001000000000000000000: n11850_o = 1'b0;
      31'b0000000000000100000000000000000: n11850_o = 1'b0;
      31'b0000000000000010000000000000000: n11850_o = 1'b0;
      31'b0000000000000001000000000000000: n11850_o = 1'b0;
      31'b0000000000000000100000000000000: n11850_o = 1'b0;
      31'b0000000000000000010000000000000: n11850_o = 1'b0;
      31'b0000000000000000001000000000000: n11850_o = 1'b0;
      31'b0000000000000000000100000000000: n11850_o = 1'b0;
      31'b0000000000000000000010000000000: n11850_o = 1'b0;
      31'b0000000000000000000001000000000: n11850_o = 1'b0;
      31'b0000000000000000000000100000000: n11850_o = 1'b0;
      31'b0000000000000000000000010000000: n11850_o = 1'b0;
      31'b0000000000000000000000001000000: n11850_o = 1'b0;
      31'b0000000000000000000000000100000: n11850_o = 1'b0;
      31'b0000000000000000000000000010000: n11850_o = 1'b0;
      31'b0000000000000000000000000001000: n11850_o = 1'b0;
      31'b0000000000000000000000000000100: n11850_o = 1'b0;
      31'b0000000000000000000000000000010: n11850_o = 1'b0;
      31'b0000000000000000000000000000001: n11850_o = 1'b0;
      default: n11850_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11851_o = 1'b0;
      31'b0100000000000000000000000000000: n11851_o = 1'b0;
      31'b0010000000000000000000000000000: n11851_o = 1'b0;
      31'b0001000000000000000000000000000: n11851_o = 1'b0;
      31'b0000100000000000000000000000000: n11851_o = 1'b0;
      31'b0000010000000000000000000000000: n11851_o = 1'b0;
      31'b0000001000000000000000000000000: n11851_o = 1'b0;
      31'b0000000100000000000000000000000: n11851_o = 1'b0;
      31'b0000000010000000000000000000000: n11851_o = 1'b0;
      31'b0000000001000000000000000000000: n11851_o = 1'b0;
      31'b0000000000100000000000000000000: n11851_o = n11546_o;
      31'b0000000000010000000000000000000: n11851_o = 1'b0;
      31'b0000000000001000000000000000000: n11851_o = 1'b0;
      31'b0000000000000100000000000000000: n11851_o = 1'b0;
      31'b0000000000000010000000000000000: n11851_o = 1'b0;
      31'b0000000000000001000000000000000: n11851_o = 1'b0;
      31'b0000000000000000100000000000000: n11851_o = 1'b0;
      31'b0000000000000000010000000000000: n11851_o = 1'b0;
      31'b0000000000000000001000000000000: n11851_o = 1'b0;
      31'b0000000000000000000100000000000: n11851_o = 1'b0;
      31'b0000000000000000000010000000000: n11851_o = 1'b0;
      31'b0000000000000000000001000000000: n11851_o = 1'b0;
      31'b0000000000000000000000100000000: n11851_o = 1'b0;
      31'b0000000000000000000000010000000: n11851_o = 1'b0;
      31'b0000000000000000000000001000000: n11851_o = 1'b0;
      31'b0000000000000000000000000100000: n11851_o = 1'b0;
      31'b0000000000000000000000000010000: n11851_o = 1'b0;
      31'b0000000000000000000000000001000: n11851_o = 1'b0;
      31'b0000000000000000000000000000100: n11851_o = 1'b0;
      31'b0000000000000000000000000000010: n11851_o = 1'b0;
      31'b0000000000000000000000000000001: n11851_o = 1'b0;
      default: n11851_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11852_o = 1'b0;
      31'b0100000000000000000000000000000: n11852_o = 1'b0;
      31'b0010000000000000000000000000000: n11852_o = 1'b0;
      31'b0001000000000000000000000000000: n11852_o = 1'b0;
      31'b0000100000000000000000000000000: n11852_o = 1'b0;
      31'b0000010000000000000000000000000: n11852_o = 1'b0;
      31'b0000001000000000000000000000000: n11852_o = n11730_o;
      31'b0000000100000000000000000000000: n11852_o = 1'b0;
      31'b0000000010000000000000000000000: n11852_o = 1'b0;
      31'b0000000001000000000000000000000: n11852_o = 1'b0;
      31'b0000000000100000000000000000000: n11852_o = 1'b0;
      31'b0000000000010000000000000000000: n11852_o = 1'b0;
      31'b0000000000001000000000000000000: n11852_o = 1'b0;
      31'b0000000000000100000000000000000: n11852_o = 1'b0;
      31'b0000000000000010000000000000000: n11852_o = 1'b0;
      31'b0000000000000001000000000000000: n11852_o = 1'b0;
      31'b0000000000000000100000000000000: n11852_o = 1'b0;
      31'b0000000000000000010000000000000: n11852_o = 1'b0;
      31'b0000000000000000001000000000000: n11852_o = 1'b0;
      31'b0000000000000000000100000000000: n11852_o = 1'b0;
      31'b0000000000000000000010000000000: n11852_o = 1'b0;
      31'b0000000000000000000001000000000: n11852_o = 1'b0;
      31'b0000000000000000000000100000000: n11852_o = 1'b0;
      31'b0000000000000000000000010000000: n11852_o = 1'b0;
      31'b0000000000000000000000001000000: n11852_o = 1'b0;
      31'b0000000000000000000000000100000: n11852_o = 1'b0;
      31'b0000000000000000000000000010000: n11852_o = 1'b0;
      31'b0000000000000000000000000001000: n11852_o = 1'b0;
      31'b0000000000000000000000000000100: n11852_o = 1'b0;
      31'b0000000000000000000000000000010: n11852_o = 1'b0;
      31'b0000000000000000000000000000001: n11852_o = 1'b0;
      default: n11852_o = 1'b0;
    endcase
  assign n11853_o = n11175_o[0];
  assign n11854_o = n11747_o[0];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11855_o = 1'b0;
      31'b0100000000000000000000000000000: n11855_o = 1'b0;
      31'b0010000000000000000000000000000: n11855_o = 1'b1;
      31'b0001000000000000000000000000000: n11855_o = 1'b1;
      31'b0000100000000000000000000000000: n11855_o = 1'b1;
      31'b0000010000000000000000000000000: n11855_o = n11854_o;
      31'b0000001000000000000000000000000: n11855_o = 1'b1;
      31'b0000000100000000000000000000000: n11855_o = 1'b1;
      31'b0000000010000000000000000000000: n11855_o = 1'b1;
      31'b0000000001000000000000000000000: n11855_o = 1'b1;
      31'b0000000000100000000000000000000: n11855_o = 1'b1;
      31'b0000000000010000000000000000000: n11855_o = 1'b1;
      31'b0000000000001000000000000000000: n11855_o = 1'b1;
      31'b0000000000000100000000000000000: n11855_o = 1'b1;
      31'b0000000000000010000000000000000: n11855_o = 1'b1;
      31'b0000000000000001000000000000000: n11855_o = 1'b1;
      31'b0000000000000000100000000000000: n11855_o = 1'b0;
      31'b0000000000000000010000000000000: n11855_o = 1'b1;
      31'b0000000000000000001000000000000: n11855_o = 1'b1;
      31'b0000000000000000000100000000000: n11855_o = 1'b1;
      31'b0000000000000000000010000000000: n11855_o = 1'b1;
      31'b0000000000000000000001000000000: n11855_o = 1'b1;
      31'b0000000000000000000000100000000: n11855_o = 1'b1;
      31'b0000000000000000000000010000000: n11855_o = 1'b1;
      31'b0000000000000000000000001000000: n11855_o = 1'b1;
      31'b0000000000000000000000000100000: n11855_o = 1'b1;
      31'b0000000000000000000000000010000: n11855_o = n11853_o;
      31'b0000000000000000000000000001000: n11855_o = 1'b1;
      31'b0000000000000000000000000000100: n11855_o = 1'b1;
      31'b0000000000000000000000000000010: n11855_o = 1'b1;
      31'b0000000000000000000000000000001: n11855_o = 1'b1;
      default: n11855_o = 1'b1;
    endcase
  assign n11856_o = n11175_o[119:1];
  assign n11857_o = n11747_o[119:1];
  assign n11858_o = {n10826_o, n10825_o, n10829_o, n10828_o};
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11859_o = n11858_o;
      31'b0100000000000000000000000000000: n11859_o = n11858_o;
      31'b0010000000000000000000000000000: n11859_o = n11858_o;
      31'b0001000000000000000000000000000: n11859_o = n11858_o;
      31'b0000100000000000000000000000000: n11859_o = n11858_o;
      31'b0000010000000000000000000000000: n11859_o = n11857_o;
      31'b0000001000000000000000000000000: n11859_o = n11858_o;
      31'b0000000100000000000000000000000: n11859_o = n11858_o;
      31'b0000000010000000000000000000000: n11859_o = n11858_o;
      31'b0000000001000000000000000000000: n11859_o = n11858_o;
      31'b0000000000100000000000000000000: n11859_o = n11858_o;
      31'b0000000000010000000000000000000: n11859_o = n11858_o;
      31'b0000000000001000000000000000000: n11859_o = n11858_o;
      31'b0000000000000100000000000000000: n11859_o = n11858_o;
      31'b0000000000000010000000000000000: n11859_o = n11858_o;
      31'b0000000000000001000000000000000: n11859_o = n11858_o;
      31'b0000000000000000100000000000000: n11859_o = n11858_o;
      31'b0000000000000000010000000000000: n11859_o = n11858_o;
      31'b0000000000000000001000000000000: n11859_o = n11858_o;
      31'b0000000000000000000100000000000: n11859_o = n11858_o;
      31'b0000000000000000000010000000000: n11859_o = n11858_o;
      31'b0000000000000000000001000000000: n11859_o = n11858_o;
      31'b0000000000000000000000100000000: n11859_o = n11858_o;
      31'b0000000000000000000000010000000: n11859_o = n11858_o;
      31'b0000000000000000000000001000000: n11859_o = n11858_o;
      31'b0000000000000000000000000100000: n11859_o = n11858_o;
      31'b0000000000000000000000000010000: n11859_o = n11856_o;
      31'b0000000000000000000000000001000: n11859_o = n11858_o;
      31'b0000000000000000000000000000100: n11859_o = n11858_o;
      31'b0000000000000000000000000000010: n11859_o = n11858_o;
      31'b0000000000000000000000000000001: n11859_o = n11858_o;
      default: n11859_o = n11858_o;
    endcase
  assign n11860_o = n11175_o[124:120];
  assign n11861_o = n11747_o[124:120];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11862_o = xerc_in;
      31'b0100000000000000000000000000000: n11862_o = xerc_in;
      31'b0010000000000000000000000000000: n11862_o = xerc_in;
      31'b0001000000000000000000000000000: n11862_o = xerc_in;
      31'b0000100000000000000000000000000: n11862_o = xerc_in;
      31'b0000010000000000000000000000000: n11862_o = n11861_o;
      31'b0000001000000000000000000000000: n11862_o = n11637_o;
      31'b0000000100000000000000000000000: n11862_o = xerc_in;
      31'b0000000010000000000000000000000: n11862_o = xerc_in;
      31'b0000000001000000000000000000000: n11862_o = xerc_in;
      31'b0000000000100000000000000000000: n11862_o = xerc_in;
      31'b0000000000010000000000000000000: n11862_o = xerc_in;
      31'b0000000000001000000000000000000: n11862_o = xerc_in;
      31'b0000000000000100000000000000000: n11862_o = xerc_in;
      31'b0000000000000010000000000000000: n11862_o = xerc_in;
      31'b0000000000000001000000000000000: n11862_o = xerc_in;
      31'b0000000000000000100000000000000: n11862_o = xerc_in;
      31'b0000000000000000010000000000000: n11862_o = xerc_in;
      31'b0000000000000000001000000000000: n11862_o = xerc_in;
      31'b0000000000000000000100000000000: n11862_o = xerc_in;
      31'b0000000000000000000010000000000: n11862_o = xerc_in;
      31'b0000000000000000000001000000000: n11862_o = xerc_in;
      31'b0000000000000000000000100000000: n11862_o = xerc_in;
      31'b0000000000000000000000010000000: n11862_o = xerc_in;
      31'b0000000000000000000000001000000: n11862_o = xerc_in;
      31'b0000000000000000000000000100000: n11862_o = xerc_in;
      31'b0000000000000000000000000010000: n11862_o = n11860_o;
      31'b0000000000000000000000000001000: n11862_o = xerc_in;
      31'b0000000000000000000000000000100: n11862_o = xerc_in;
      31'b0000000000000000000000000000010: n11862_o = xerc_in;
      31'b0000000000000000000000000000001: n11862_o = xerc_in;
      default: n11862_o = xerc_in;
    endcase
  assign n11863_o = n11175_o[125];
  assign n11864_o = n11747_o[125];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11865_o = n10816_o;
      31'b0100000000000000000000000000000: n11865_o = n10816_o;
      31'b0010000000000000000000000000000: n11865_o = n10816_o;
      31'b0001000000000000000000000000000: n11865_o = n10816_o;
      31'b0000100000000000000000000000000: n11865_o = n10816_o;
      31'b0000010000000000000000000000000: n11865_o = n11864_o;
      31'b0000001000000000000000000000000: n11865_o = n10816_o;
      31'b0000000100000000000000000000000: n11865_o = n10816_o;
      31'b0000000010000000000000000000000: n11865_o = n10816_o;
      31'b0000000001000000000000000000000: n11865_o = n10816_o;
      31'b0000000000100000000000000000000: n11865_o = n10816_o;
      31'b0000000000010000000000000000000: n11865_o = n10816_o;
      31'b0000000000001000000000000000000: n11865_o = n10816_o;
      31'b0000000000000100000000000000000: n11865_o = n10816_o;
      31'b0000000000000010000000000000000: n11865_o = n10816_o;
      31'b0000000000000001000000000000000: n11865_o = n10816_o;
      31'b0000000000000000100000000000000: n11865_o = n10816_o;
      31'b0000000000000000010000000000000: n11865_o = n10816_o;
      31'b0000000000000000001000000000000: n11865_o = n10816_o;
      31'b0000000000000000000100000000000: n11865_o = n10816_o;
      31'b0000000000000000000010000000000: n11865_o = n10816_o;
      31'b0000000000000000000001000000000: n11865_o = n10816_o;
      31'b0000000000000000000000100000000: n11865_o = n10816_o;
      31'b0000000000000000000000010000000: n11865_o = n10816_o;
      31'b0000000000000000000000001000000: n11865_o = n10816_o;
      31'b0000000000000000000000000100000: n11865_o = n10816_o;
      31'b0000000000000000000000000010000: n11865_o = n11863_o;
      31'b0000000000000000000000000001000: n11865_o = n10816_o;
      31'b0000000000000000000000000000100: n11865_o = n10816_o;
      31'b0000000000000000000000000000010: n11865_o = n10816_o;
      31'b0000000000000000000000000000001: n11865_o = n10816_o;
      default: n11865_o = n10816_o;
    endcase
  assign n11866_o = n11175_o[137:126];
  assign n11867_o = n11747_o[137:126];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11868_o = n11011_o;
      31'b0100000000000000000000000000000: n11868_o = n11011_o;
      31'b0010000000000000000000000000000: n11868_o = n11011_o;
      31'b0001000000000000000000000000000: n11868_o = n11011_o;
      31'b0000100000000000000000000000000: n11868_o = n11011_o;
      31'b0000010000000000000000000000000: n11868_o = n11867_o;
      31'b0000001000000000000000000000000: n11868_o = n11011_o;
      31'b0000000100000000000000000000000: n11868_o = n11011_o;
      31'b0000000010000000000000000000000: n11868_o = n11011_o;
      31'b0000000001000000000000000000000: n11868_o = n11011_o;
      31'b0000000000100000000000000000000: n11868_o = n11011_o;
      31'b0000000000010000000000000000000: n11868_o = n11011_o;
      31'b0000000000001000000000000000000: n11868_o = n11011_o;
      31'b0000000000000100000000000000000: n11868_o = n11011_o;
      31'b0000000000000010000000000000000: n11868_o = n11011_o;
      31'b0000000000000001000000000000000: n11868_o = n11011_o;
      31'b0000000000000000100000000000000: n11868_o = n11011_o;
      31'b0000000000000000010000000000000: n11868_o = n11011_o;
      31'b0000000000000000001000000000000: n11868_o = n11011_o;
      31'b0000000000000000000100000000000: n11868_o = n11011_o;
      31'b0000000000000000000010000000000: n11868_o = n11011_o;
      31'b0000000000000000000001000000000: n11868_o = n11011_o;
      31'b0000000000000000000000100000000: n11868_o = n11011_o;
      31'b0000000000000000000000010000000: n11868_o = n11011_o;
      31'b0000000000000000000000001000000: n11868_o = 12'b011100000000;
      31'b0000000000000000000000000100000: n11868_o = n11011_o;
      31'b0000000000000000000000000010000: n11868_o = n11866_o;
      31'b0000000000000000000000000001000: n11868_o = n11011_o;
      31'b0000000000000000000000000000100: n11868_o = n11011_o;
      31'b0000000000000000000000000000010: n11868_o = n11101_o;
      31'b0000000000000000000000000000001: n11868_o = n11011_o;
      default: n11868_o = n11011_o;
    endcase
  assign n11869_o = n11175_o[138];
  assign n11870_o = n11747_o[138];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11871_o = n10815_o;
      31'b0100000000000000000000000000000: n11871_o = n10815_o;
      31'b0010000000000000000000000000000: n11871_o = n10815_o;
      31'b0001000000000000000000000000000: n11871_o = 1'b1;
      31'b0000100000000000000000000000000: n11871_o = n10815_o;
      31'b0000010000000000000000000000000: n11871_o = n11870_o;
      31'b0000001000000000000000000000000: n11871_o = n10815_o;
      31'b0000000100000000000000000000000: n11871_o = n10815_o;
      31'b0000000010000000000000000000000: n11871_o = n10815_o;
      31'b0000000001000000000000000000000: n11871_o = n10815_o;
      31'b0000000000100000000000000000000: n11871_o = n10815_o;
      31'b0000000000010000000000000000000: n11871_o = n10815_o;
      31'b0000000000001000000000000000000: n11871_o = n10815_o;
      31'b0000000000000100000000000000000: n11871_o = n10815_o;
      31'b0000000000000010000000000000000: n11871_o = n10815_o;
      31'b0000000000000001000000000000000: n11871_o = n10815_o;
      31'b0000000000000000100000000000000: n11871_o = n10815_o;
      31'b0000000000000000010000000000000: n11871_o = n10815_o;
      31'b0000000000000000001000000000000: n11871_o = n10815_o;
      31'b0000000000000000000100000000000: n11871_o = n10815_o;
      31'b0000000000000000000010000000000: n11871_o = n10815_o;
      31'b0000000000000000000001000000000: n11871_o = n10815_o;
      31'b0000000000000000000000100000000: n11871_o = n10815_o;
      31'b0000000000000000000000010000000: n11871_o = n10815_o;
      31'b0000000000000000000000001000000: n11871_o = n10815_o;
      31'b0000000000000000000000000100000: n11871_o = n10815_o;
      31'b0000000000000000000000000010000: n11871_o = n11869_o;
      31'b0000000000000000000000000001000: n11871_o = n10815_o;
      31'b0000000000000000000000000000100: n11871_o = n10815_o;
      31'b0000000000000000000000000000010: n11871_o = n10815_o;
      31'b0000000000000000000000000000001: n11871_o = n10815_o;
      default: n11871_o = n10815_o;
    endcase
  assign n11872_o = n11175_o[142:139];
  assign n11873_o = n11747_o[142:139];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11874_o = n10715_o;
      31'b0100000000000000000000000000000: n11874_o = n10715_o;
      31'b0010000000000000000000000000000: n11874_o = n10715_o;
      31'b0001000000000000000000000000000: n11874_o = n10715_o;
      31'b0000100000000000000000000000000: n11874_o = n10715_o;
      31'b0000010000000000000000000000000: n11874_o = n11873_o;
      31'b0000001000000000000000000000000: n11874_o = n10715_o;
      31'b0000000100000000000000000000000: n11874_o = n10715_o;
      31'b0000000010000000000000000000000: n11874_o = n10715_o;
      31'b0000000001000000000000000000000: n11874_o = n10715_o;
      31'b0000000000100000000000000000000: n11874_o = n10715_o;
      31'b0000000000010000000000000000000: n11874_o = n10715_o;
      31'b0000000000001000000000000000000: n11874_o = n10715_o;
      31'b0000000000000100000000000000000: n11874_o = n10715_o;
      31'b0000000000000010000000000000000: n11874_o = n10715_o;
      31'b0000000000000001000000000000000: n11874_o = n10715_o;
      31'b0000000000000000100000000000000: n11874_o = n10715_o;
      31'b0000000000000000010000000000000: n11874_o = n11324_o;
      31'b0000000000000000001000000000000: n11874_o = n10715_o;
      31'b0000000000000000000100000000000: n11874_o = n10715_o;
      31'b0000000000000000000010000000000: n11874_o = n10715_o;
      31'b0000000000000000000001000000000: n11874_o = n10715_o;
      31'b0000000000000000000000100000000: n11874_o = n10715_o;
      31'b0000000000000000000000010000000: n11874_o = n10715_o;
      31'b0000000000000000000000001000000: n11874_o = n10715_o;
      31'b0000000000000000000000000100000: n11874_o = n10715_o;
      31'b0000000000000000000000000010000: n11874_o = n11872_o;
      31'b0000000000000000000000000001000: n11874_o = n10715_o;
      31'b0000000000000000000000000000100: n11874_o = n10715_o;
      31'b0000000000000000000000000000010: n11874_o = n10715_o;
      31'b0000000000000000000000000000001: n11874_o = n10715_o;
      default: n11874_o = n10715_o;
    endcase
  assign n11875_o = n11175_o[206:143];
  assign n11876_o = n11747_o[206:143];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11877_o = n10822_o;
      31'b0100000000000000000000000000000: n11877_o = n10822_o;
      31'b0010000000000000000000000000000: n11877_o = n10822_o;
      31'b0001000000000000000000000000000: n11877_o = n10822_o;
      31'b0000100000000000000000000000000: n11877_o = n10822_o;
      31'b0000010000000000000000000000000: n11877_o = n11876_o;
      31'b0000001000000000000000000000000: n11877_o = n10822_o;
      31'b0000000100000000000000000000000: n11877_o = n10822_o;
      31'b0000000010000000000000000000000: n11877_o = n10822_o;
      31'b0000000001000000000000000000000: n11877_o = n10822_o;
      31'b0000000000100000000000000000000: n11877_o = n10822_o;
      31'b0000000000010000000000000000000: n11877_o = n10822_o;
      31'b0000000000001000000000000000000: n11877_o = n10822_o;
      31'b0000000000000100000000000000000: n11877_o = n10822_o;
      31'b0000000000000010000000000000000: n11877_o = n10822_o;
      31'b0000000000000001000000000000000: n11877_o = n10822_o;
      31'b0000000000000000100000000000000: n11877_o = n10822_o;
      31'b0000000000000000010000000000000: n11877_o = n10822_o;
      31'b0000000000000000001000000000000: n11877_o = n10822_o;
      31'b0000000000000000000100000000000: n11877_o = n10822_o;
      31'b0000000000000000000010000000000: n11877_o = n10822_o;
      31'b0000000000000000000001000000000: n11877_o = n10822_o;
      31'b0000000000000000000000100000000: n11877_o = n10822_o;
      31'b0000000000000000000000010000000: n11877_o = n10822_o;
      31'b0000000000000000000000001000000: n11877_o = n10822_o;
      31'b0000000000000000000000000100000: n11877_o = n10822_o;
      31'b0000000000000000000000000010000: n11877_o = n11875_o;
      31'b0000000000000000000000000001000: n11877_o = n10822_o;
      31'b0000000000000000000000000000100: n11877_o = n10822_o;
      31'b0000000000000000000000000000010: n11877_o = n11102_o;
      31'b0000000000000000000000000000001: n11877_o = n10822_o;
      default: n11877_o = n10822_o;
    endcase
  assign n11878_o = n11175_o[270:207];
  assign n11879_o = n11747_o[270:207];
  assign n11880_o = n10704_o[270:207];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11881_o = n11880_o;
      31'b0100000000000000000000000000000: n11881_o = n11880_o;
      31'b0010000000000000000000000000000: n11881_o = n11880_o;
      31'b0001000000000000000000000000000: n11881_o = 64'b0000000000000000000000000000000000000000000000000000000000000100;
      31'b0000100000000000000000000000000: n11881_o = n11880_o;
      31'b0000010000000000000000000000000: n11881_o = n11879_o;
      31'b0000001000000000000000000000000: n11881_o = n11880_o;
      31'b0000000100000000000000000000000: n11881_o = n11880_o;
      31'b0000000010000000000000000000000: n11881_o = n11880_o;
      31'b0000000001000000000000000000000: n11881_o = n11880_o;
      31'b0000000000100000000000000000000: n11881_o = n11880_o;
      31'b0000000000010000000000000000000: n11881_o = n11880_o;
      31'b0000000000001000000000000000000: n11881_o = n11880_o;
      31'b0000000000000100000000000000000: n11881_o = n11880_o;
      31'b0000000000000010000000000000000: n11881_o = n11880_o;
      31'b0000000000000001000000000000000: n11881_o = n11880_o;
      31'b0000000000000000100000000000000: n11881_o = n11880_o;
      31'b0000000000000000010000000000000: n11881_o = n11880_o;
      31'b0000000000000000001000000000000: n11881_o = n11880_o;
      31'b0000000000000000000100000000000: n11881_o = n11880_o;
      31'b0000000000000000000010000000000: n11881_o = n11880_o;
      31'b0000000000000000000001000000000: n11881_o = n11880_o;
      31'b0000000000000000000000100000000: n11881_o = n11880_o;
      31'b0000000000000000000000010000000: n11881_o = n11880_o;
      31'b0000000000000000000000001000000: n11881_o = n11880_o;
      31'b0000000000000000000000000100000: n11881_o = n11880_o;
      31'b0000000000000000000000000010000: n11881_o = n11878_o;
      31'b0000000000000000000000000001000: n11881_o = n11880_o;
      31'b0000000000000000000000000000100: n11881_o = n11880_o;
      31'b0000000000000000000000000000010: n11881_o = n11880_o;
      31'b0000000000000000000000000000001: n11881_o = n11880_o;
      default: n11881_o = n11880_o;
    endcase
  assign n11882_o = n11175_o[274:271];
  assign n11883_o = n11747_o[274:271];
  assign n11884_o = n10704_o[273:271];
  assign n11885_o = {n11015_o, n11884_o};
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11886_o = n11885_o;
      31'b0100000000000000000000000000000: n11886_o = n11885_o;
      31'b0010000000000000000000000000000: n11886_o = n11885_o;
      31'b0001000000000000000000000000000: n11886_o = n11885_o;
      31'b0000100000000000000000000000000: n11886_o = n11885_o;
      31'b0000010000000000000000000000000: n11886_o = n11883_o;
      31'b0000001000000000000000000000000: n11886_o = n11885_o;
      31'b0000000100000000000000000000000: n11886_o = n11885_o;
      31'b0000000010000000000000000000000: n11886_o = n11885_o;
      31'b0000000001000000000000000000000: n11886_o = n11885_o;
      31'b0000000000100000000000000000000: n11886_o = n11885_o;
      31'b0000000000010000000000000000000: n11886_o = n11885_o;
      31'b0000000000001000000000000000000: n11886_o = n11885_o;
      31'b0000000000000100000000000000000: n11886_o = n11885_o;
      31'b0000000000000010000000000000000: n11886_o = n11885_o;
      31'b0000000000000001000000000000000: n11886_o = n11885_o;
      31'b0000000000000000100000000000000: n11886_o = n11885_o;
      31'b0000000000000000010000000000000: n11886_o = n11885_o;
      31'b0000000000000000001000000000000: n11886_o = n11885_o;
      31'b0000000000000000000100000000000: n11886_o = n11885_o;
      31'b0000000000000000000010000000000: n11886_o = n11885_o;
      31'b0000000000000000000001000000000: n11886_o = n11885_o;
      31'b0000000000000000000000100000000: n11886_o = n11885_o;
      31'b0000000000000000000000010000000: n11886_o = n11885_o;
      31'b0000000000000000000000001000000: n11886_o = n11885_o;
      31'b0000000000000000000000000100000: n11886_o = n11885_o;
      31'b0000000000000000000000000010000: n11886_o = n11882_o;
      31'b0000000000000000000000000001000: n11886_o = n11885_o;
      31'b0000000000000000000000000000100: n11886_o = n11885_o;
      31'b0000000000000000000000000000010: n11886_o = n11885_o;
      31'b0000000000000000000000000000001: n11886_o = n11885_o;
      default: n11886_o = n11885_o;
    endcase
  assign n11887_o = n11175_o[275];
  assign n11888_o = n11747_o[275];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11889_o = n11041_o;
      31'b0100000000000000000000000000000: n11889_o = n11041_o;
      31'b0010000000000000000000000000000: n11889_o = n11041_o;
      31'b0001000000000000000000000000000: n11889_o = n11041_o;
      31'b0000100000000000000000000000000: n11889_o = n11041_o;
      31'b0000010000000000000000000000000: n11889_o = n11888_o;
      31'b0000001000000000000000000000000: n11889_o = n11041_o;
      31'b0000000100000000000000000000000: n11889_o = n11041_o;
      31'b0000000010000000000000000000000: n11889_o = n11041_o;
      31'b0000000001000000000000000000000: n11889_o = n11041_o;
      31'b0000000000100000000000000000000: n11889_o = n11041_o;
      31'b0000000000010000000000000000000: n11889_o = n11041_o;
      31'b0000000000001000000000000000000: n11889_o = n11041_o;
      31'b0000000000000100000000000000000: n11889_o = n11041_o;
      31'b0000000000000010000000000000000: n11889_o = n11041_o;
      31'b0000000000000001000000000000000: n11889_o = n11041_o;
      31'b0000000000000000100000000000000: n11889_o = n11041_o;
      31'b0000000000000000010000000000000: n11889_o = n11041_o;
      31'b0000000000000000001000000000000: n11889_o = n11041_o;
      31'b0000000000000000000100000000000: n11889_o = n11041_o;
      31'b0000000000000000000010000000000: n11889_o = n11041_o;
      31'b0000000000000000000001000000000: n11889_o = n11041_o;
      31'b0000000000000000000000100000000: n11889_o = n11041_o;
      31'b0000000000000000000000010000000: n11889_o = n11041_o;
      31'b0000000000000000000000001000000: n11889_o = 1'b1;
      31'b0000000000000000000000000100000: n11889_o = n11041_o;
      31'b0000000000000000000000000010000: n11889_o = n11887_o;
      31'b0000000000000000000000000001000: n11889_o = n11041_o;
      31'b0000000000000000000000000000100: n11889_o = n11041_o;
      31'b0000000000000000000000000000010: n11889_o = n11041_o;
      31'b0000000000000000000000000000001: n11889_o = n11041_o;
      default: n11889_o = n11041_o;
    endcase
  assign n11890_o = n11175_o[353:276];
  assign n11891_o = n11747_o[353:276];
  assign n11892_o = {n10817_o, n11056_o, n11031_o, n11059_o, n11027_o, n11053_o, n11023_o, n11047_o, n11019_o};
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11893_o = n11892_o;
      31'b0100000000000000000000000000000: n11893_o = n11892_o;
      31'b0010000000000000000000000000000: n11893_o = n11892_o;
      31'b0001000000000000000000000000000: n11893_o = n11892_o;
      31'b0000100000000000000000000000000: n11893_o = n11892_o;
      31'b0000010000000000000000000000000: n11893_o = n11891_o;
      31'b0000001000000000000000000000000: n11893_o = n11892_o;
      31'b0000000100000000000000000000000: n11893_o = n11892_o;
      31'b0000000010000000000000000000000: n11893_o = n11892_o;
      31'b0000000001000000000000000000000: n11893_o = n11892_o;
      31'b0000000000100000000000000000000: n11893_o = n11892_o;
      31'b0000000000010000000000000000000: n11893_o = n11892_o;
      31'b0000000000001000000000000000000: n11893_o = n11892_o;
      31'b0000000000000100000000000000000: n11893_o = n11892_o;
      31'b0000000000000010000000000000000: n11893_o = n11892_o;
      31'b0000000000000001000000000000000: n11893_o = n11892_o;
      31'b0000000000000000100000000000000: n11893_o = n11892_o;
      31'b0000000000000000010000000000000: n11893_o = n11892_o;
      31'b0000000000000000001000000000000: n11893_o = n11892_o;
      31'b0000000000000000000100000000000: n11893_o = n11892_o;
      31'b0000000000000000000010000000000: n11893_o = n11892_o;
      31'b0000000000000000000001000000000: n11893_o = n11892_o;
      31'b0000000000000000000000100000000: n11893_o = n11892_o;
      31'b0000000000000000000000010000000: n11893_o = n11892_o;
      31'b0000000000000000000000001000000: n11893_o = n11892_o;
      31'b0000000000000000000000000100000: n11893_o = n11892_o;
      31'b0000000000000000000000000010000: n11893_o = n11890_o;
      31'b0000000000000000000000000001000: n11893_o = n11892_o;
      31'b0000000000000000000000000000100: n11893_o = n11892_o;
      31'b0000000000000000000000000000010: n11893_o = n11892_o;
      31'b0000000000000000000000000000001: n11893_o = n11892_o;
      default: n11893_o = n11892_o;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11894_o = 1'b1;
      31'b0100000000000000000000000000000: n11894_o = 1'b1;
      31'b0010000000000000000000000000000: n11894_o = n11065_o;
      31'b0001000000000000000000000000000: n11894_o = n11065_o;
      31'b0000100000000000000000000000000: n11894_o = n11065_o;
      31'b0000010000000000000000000000000: n11894_o = n11065_o;
      31'b0000001000000000000000000000000: n11894_o = n11065_o;
      31'b0000000100000000000000000000000: n11894_o = n11065_o;
      31'b0000000010000000000000000000000: n11894_o = n11065_o;
      31'b0000000001000000000000000000000: n11894_o = n11065_o;
      31'b0000000000100000000000000000000: n11894_o = n11065_o;
      31'b0000000000010000000000000000000: n11894_o = n11065_o;
      31'b0000000000001000000000000000000: n11894_o = n11065_o;
      31'b0000000000000100000000000000000: n11894_o = n11065_o;
      31'b0000000000000010000000000000000: n11894_o = n11065_o;
      31'b0000000000000001000000000000000: n11894_o = n11065_o;
      31'b0000000000000000100000000000000: n11894_o = 1'b1;
      31'b0000000000000000010000000000000: n11894_o = n11065_o;
      31'b0000000000000000001000000000000: n11894_o = n11065_o;
      31'b0000000000000000000100000000000: n11894_o = n11065_o;
      31'b0000000000000000000010000000000: n11894_o = n11065_o;
      31'b0000000000000000000001000000000: n11894_o = n11065_o;
      31'b0000000000000000000000100000000: n11894_o = n11065_o;
      31'b0000000000000000000000010000000: n11894_o = n11065_o;
      31'b0000000000000000000000001000000: n11894_o = n11065_o;
      31'b0000000000000000000000000100000: n11894_o = n11065_o;
      31'b0000000000000000000000000010000: n11894_o = n11065_o;
      31'b0000000000000000000000000001000: n11894_o = n11065_o;
      31'b0000000000000000000000000000100: n11894_o = n11065_o;
      31'b0000000000000000000000000000010: n11894_o = n11065_o;
      31'b0000000000000000000000000000001: n11894_o = n11065_o;
      default: n11894_o = n11065_o;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11895_o = 1'b0;
      31'b0100000000000000000000000000000: n11895_o = 1'b0;
      31'b0010000000000000000000000000000: n11895_o = 1'b0;
      31'b0001000000000000000000000000000: n11895_o = 1'b0;
      31'b0000100000000000000000000000000: n11895_o = 1'b0;
      31'b0000010000000000000000000000000: n11895_o = 1'b0;
      31'b0000001000000000000000000000000: n11895_o = 1'b0;
      31'b0000000100000000000000000000000: n11895_o = 1'b0;
      31'b0000000010000000000000000000000: n11895_o = 1'b0;
      31'b0000000001000000000000000000000: n11895_o = 1'b0;
      31'b0000000000100000000000000000000: n11895_o = 1'b0;
      31'b0000000000010000000000000000000: n11895_o = 1'b0;
      31'b0000000000001000000000000000000: n11895_o = 1'b0;
      31'b0000000000000100000000000000000: n11895_o = 1'b0;
      31'b0000000000000010000000000000000: n11895_o = 1'b0;
      31'b0000000000000001000000000000000: n11895_o = 1'b0;
      31'b0000000000000000100000000000000: n11895_o = 1'b0;
      31'b0000000000000000010000000000000: n11895_o = 1'b0;
      31'b0000000000000000001000000000000: n11895_o = 1'b0;
      31'b0000000000000000000100000000000: n11895_o = 1'b0;
      31'b0000000000000000000010000000000: n11895_o = 1'b0;
      31'b0000000000000000000001000000000: n11895_o = 1'b0;
      31'b0000000000000000000000100000000: n11895_o = 1'b0;
      31'b0000000000000000000000010000000: n11895_o = 1'b0;
      31'b0000000000000000000000001000000: n11895_o = 1'b0;
      31'b0000000000000000000000000100000: n11895_o = 1'b0;
      31'b0000000000000000000000000010000: n11895_o = 1'b0;
      31'b0000000000000000000000000001000: n11895_o = 1'b0;
      31'b0000000000000000000000000000100: n11895_o = n11114_o;
      31'b0000000000000000000000000000010: n11895_o = 1'b0;
      31'b0000000000000000000000000000001: n11895_o = 1'b0;
      default: n11895_o = 1'b1;
    endcase
  assign n11896_o = r[749];
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11897_o = n11896_o;
      31'b0100000000000000000000000000000: n11897_o = n11896_o;
      31'b0010000000000000000000000000000: n11897_o = n11896_o;
      31'b0001000000000000000000000000000: n11897_o = n11896_o;
      31'b0000100000000000000000000000000: n11897_o = n11896_o;
      31'b0000010000000000000000000000000: n11897_o = n11896_o;
      31'b0000001000000000000000000000000: n11897_o = n11896_o;
      31'b0000000100000000000000000000000: n11897_o = n11608_o;
      31'b0000000010000000000000000000000: n11897_o = n11896_o;
      31'b0000000001000000000000000000000: n11897_o = n11896_o;
      31'b0000000000100000000000000000000: n11897_o = n11896_o;
      31'b0000000000010000000000000000000: n11897_o = n11896_o;
      31'b0000000000001000000000000000000: n11897_o = n11896_o;
      31'b0000000000000100000000000000000: n11897_o = n11896_o;
      31'b0000000000000010000000000000000: n11897_o = n11896_o;
      31'b0000000000000001000000000000000: n11897_o = n11896_o;
      31'b0000000000000000100000000000000: n11897_o = n11896_o;
      31'b0000000000000000010000000000000: n11897_o = n11344_o;
      31'b0000000000000000001000000000000: n11897_o = n11896_o;
      31'b0000000000000000000100000000000: n11897_o = n11896_o;
      31'b0000000000000000000010000000000: n11897_o = n11896_o;
      31'b0000000000000000000001000000000: n11897_o = n11896_o;
      31'b0000000000000000000000100000000: n11897_o = n11896_o;
      31'b0000000000000000000000010000000: n11897_o = n11896_o;
      31'b0000000000000000000000001000000: n11897_o = n11896_o;
      31'b0000000000000000000000000100000: n11897_o = n11896_o;
      31'b0000000000000000000000000010000: n11897_o = n11896_o;
      31'b0000000000000000000000000001000: n11897_o = n11896_o;
      31'b0000000000000000000000000000100: n11897_o = n11896_o;
      31'b0000000000000000000000000000010: n11897_o = n11896_o;
      31'b0000000000000000000000000000001: n11897_o = n11896_o;
      default: n11897_o = n11896_o;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11898_o = n10837_o;
      31'b0100000000000000000000000000000: n11898_o = n10837_o;
      31'b0010000000000000000000000000000: n11898_o = n10837_o;
      31'b0001000000000000000000000000000: n11898_o = n10837_o;
      31'b0000100000000000000000000000000: n11898_o = n10837_o;
      31'b0000010000000000000000000000000: n11898_o = n10837_o;
      31'b0000001000000000000000000000000: n11898_o = n10837_o;
      31'b0000000100000000000000000000000: n11898_o = n10837_o;
      31'b0000000010000000000000000000000: n11898_o = n10837_o;
      31'b0000000001000000000000000000000: n11898_o = n10837_o;
      31'b0000000000100000000000000000000: n11898_o = n10837_o;
      31'b0000000000010000000000000000000: n11898_o = n10837_o;
      31'b0000000000001000000000000000000: n11898_o = n10837_o;
      31'b0000000000000100000000000000000: n11898_o = n10837_o;
      31'b0000000000000010000000000000000: n11898_o = n10837_o;
      31'b0000000000000001000000000000000: n11898_o = n10837_o;
      31'b0000000000000000100000000000000: n11898_o = n10837_o;
      31'b0000000000000000010000000000000: n11898_o = n10837_o;
      31'b0000000000000000001000000000000: n11898_o = n11287_o;
      31'b0000000000000000000100000000000: n11898_o = n10837_o;
      31'b0000000000000000000010000000000: n11898_o = n10837_o;
      31'b0000000000000000000001000000000: n11898_o = n10837_o;
      31'b0000000000000000000000100000000: n11898_o = n10837_o;
      31'b0000000000000000000000010000000: n11898_o = n10837_o;
      31'b0000000000000000000000001000000: n11898_o = n10837_o;
      31'b0000000000000000000000000100000: n11898_o = n10837_o;
      31'b0000000000000000000000000010000: n11898_o = n10837_o;
      31'b0000000000000000000000000001000: n11898_o = n10837_o;
      31'b0000000000000000000000000000100: n11898_o = n10837_o;
      31'b0000000000000000000000000000010: n11898_o = n10837_o;
      31'b0000000000000000000000000000001: n11898_o = n10837_o;
      default: n11898_o = n10837_o;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11899_o = 1'b0;
      31'b0100000000000000000000000000000: n11899_o = 1'b1;
      31'b0010000000000000000000000000000: n11899_o = 1'b0;
      31'b0001000000000000000000000000000: n11899_o = 1'b0;
      31'b0000100000000000000000000000000: n11899_o = 1'b0;
      31'b0000010000000000000000000000000: n11899_o = 1'b0;
      31'b0000001000000000000000000000000: n11899_o = 1'b0;
      31'b0000000100000000000000000000000: n11899_o = 1'b0;
      31'b0000000010000000000000000000000: n11899_o = 1'b0;
      31'b0000000001000000000000000000000: n11899_o = 1'b0;
      31'b0000000000100000000000000000000: n11899_o = 1'b0;
      31'b0000000000010000000000000000000: n11899_o = 1'b0;
      31'b0000000000001000000000000000000: n11899_o = 1'b0;
      31'b0000000000000100000000000000000: n11899_o = 1'b0;
      31'b0000000000000010000000000000000: n11899_o = 1'b0;
      31'b0000000000000001000000000000000: n11899_o = 1'b0;
      31'b0000000000000000100000000000000: n11899_o = 1'b0;
      31'b0000000000000000010000000000000: n11899_o = 1'b0;
      31'b0000000000000000001000000000000: n11899_o = 1'b0;
      31'b0000000000000000000100000000000: n11899_o = 1'b0;
      31'b0000000000000000000010000000000: n11899_o = 1'b0;
      31'b0000000000000000000001000000000: n11899_o = 1'b0;
      31'b0000000000000000000000100000000: n11899_o = 1'b0;
      31'b0000000000000000000000010000000: n11899_o = 1'b0;
      31'b0000000000000000000000001000000: n11899_o = 1'b0;
      31'b0000000000000000000000000100000: n11899_o = 1'b0;
      31'b0000000000000000000000000010000: n11899_o = 1'b0;
      31'b0000000000000000000000000001000: n11899_o = 1'b0;
      31'b0000000000000000000000000000100: n11899_o = 1'b0;
      31'b0000000000000000000000000000010: n11899_o = 1'b0;
      31'b0000000000000000000000000000001: n11899_o = 1'b0;
      default: n11899_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11900_o = 1'b1;
      31'b0100000000000000000000000000000: n11900_o = 1'b0;
      31'b0010000000000000000000000000000: n11900_o = 1'b0;
      31'b0001000000000000000000000000000: n11900_o = 1'b0;
      31'b0000100000000000000000000000000: n11900_o = 1'b0;
      31'b0000010000000000000000000000000: n11900_o = 1'b0;
      31'b0000001000000000000000000000000: n11900_o = 1'b0;
      31'b0000000100000000000000000000000: n11900_o = 1'b0;
      31'b0000000010000000000000000000000: n11900_o = 1'b0;
      31'b0000000001000000000000000000000: n11900_o = 1'b0;
      31'b0000000000100000000000000000000: n11900_o = 1'b0;
      31'b0000000000010000000000000000000: n11900_o = 1'b0;
      31'b0000000000001000000000000000000: n11900_o = 1'b0;
      31'b0000000000000100000000000000000: n11900_o = 1'b0;
      31'b0000000000000010000000000000000: n11900_o = 1'b0;
      31'b0000000000000001000000000000000: n11900_o = 1'b0;
      31'b0000000000000000100000000000000: n11900_o = 1'b0;
      31'b0000000000000000010000000000000: n11900_o = 1'b0;
      31'b0000000000000000001000000000000: n11900_o = 1'b0;
      31'b0000000000000000000100000000000: n11900_o = 1'b0;
      31'b0000000000000000000010000000000: n11900_o = 1'b0;
      31'b0000000000000000000001000000000: n11900_o = 1'b0;
      31'b0000000000000000000000100000000: n11900_o = 1'b0;
      31'b0000000000000000000000010000000: n11900_o = 1'b0;
      31'b0000000000000000000000001000000: n11900_o = 1'b0;
      31'b0000000000000000000000000100000: n11900_o = 1'b0;
      31'b0000000000000000000000000010000: n11900_o = 1'b0;
      31'b0000000000000000000000000001000: n11900_o = 1'b0;
      31'b0000000000000000000000000000100: n11900_o = 1'b0;
      31'b0000000000000000000000000000010: n11900_o = 1'b0;
      31'b0000000000000000000000000000001: n11900_o = 1'b0;
      default: n11900_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11901_o = 1'b0;
      31'b0100000000000000000000000000000: n11901_o = 1'b0;
      31'b0010000000000000000000000000000: n11901_o = 1'b0;
      31'b0001000000000000000000000000000: n11901_o = 1'b0;
      31'b0000100000000000000000000000000: n11901_o = 1'b0;
      31'b0000010000000000000000000000000: n11901_o = 1'b0;
      31'b0000001000000000000000000000000: n11901_o = 1'b0;
      31'b0000000100000000000000000000000: n11901_o = 1'b0;
      31'b0000000010000000000000000000000: n11901_o = 1'b0;
      31'b0000000001000000000000000000000: n11901_o = 1'b0;
      31'b0000000000100000000000000000000: n11901_o = 1'b0;
      31'b0000000000010000000000000000000: n11901_o = 1'b0;
      31'b0000000000001000000000000000000: n11901_o = 1'b0;
      31'b0000000000000100000000000000000: n11901_o = 1'b0;
      31'b0000000000000010000000000000000: n11901_o = 1'b0;
      31'b0000000000000001000000000000000: n11901_o = 1'b0;
      31'b0000000000000000100000000000000: n11901_o = 1'b1;
      31'b0000000000000000010000000000000: n11901_o = 1'b0;
      31'b0000000000000000001000000000000: n11901_o = 1'b0;
      31'b0000000000000000000100000000000: n11901_o = 1'b0;
      31'b0000000000000000000010000000000: n11901_o = 1'b0;
      31'b0000000000000000000001000000000: n11901_o = 1'b0;
      31'b0000000000000000000000100000000: n11901_o = 1'b0;
      31'b0000000000000000000000010000000: n11901_o = 1'b0;
      31'b0000000000000000000000001000000: n11901_o = 1'b0;
      31'b0000000000000000000000000100000: n11901_o = 1'b0;
      31'b0000000000000000000000000010000: n11901_o = 1'b0;
      31'b0000000000000000000000000001000: n11901_o = 1'b0;
      31'b0000000000000000000000000000100: n11901_o = 1'b0;
      31'b0000000000000000000000000000010: n11901_o = 1'b0;
      31'b0000000000000000000000000000001: n11901_o = 1'b0;
      default: n11901_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11902_o = 1'b0;
      31'b0100000000000000000000000000000: n11902_o = 1'b0;
      31'b0010000000000000000000000000000: n11902_o = 1'b0;
      31'b0001000000000000000000000000000: n11902_o = 1'b0;
      31'b0000100000000000000000000000000: n11902_o = 1'b0;
      31'b0000010000000000000000000000000: n11902_o = 1'b0;
      31'b0000001000000000000000000000000: n11902_o = 1'b0;
      31'b0000000100000000000000000000000: n11902_o = 1'b0;
      31'b0000000010000000000000000000000: n11902_o = 1'b0;
      31'b0000000001000000000000000000000: n11902_o = 1'b0;
      31'b0000000000100000000000000000000: n11902_o = 1'b0;
      31'b0000000000010000000000000000000: n11902_o = 1'b0;
      31'b0000000000001000000000000000000: n11902_o = 1'b0;
      31'b0000000000000100000000000000000: n11902_o = 1'b0;
      31'b0000000000000010000000000000000: n11902_o = 1'b0;
      31'b0000000000000001000000000000000: n11902_o = 1'b0;
      31'b0000000000000000100000000000000: n11902_o = 1'b0;
      31'b0000000000000000010000000000000: n11902_o = 1'b0;
      31'b0000000000000000001000000000000: n11902_o = n11287_o;
      31'b0000000000000000000100000000000: n11902_o = 1'b1;
      31'b0000000000000000000010000000000: n11902_o = 1'b0;
      31'b0000000000000000000001000000000: n11902_o = 1'b0;
      31'b0000000000000000000000100000000: n11902_o = 1'b0;
      31'b0000000000000000000000010000000: n11902_o = 1'b0;
      31'b0000000000000000000000001000000: n11902_o = 1'b0;
      31'b0000000000000000000000000100000: n11902_o = 1'b0;
      31'b0000000000000000000000000010000: n11902_o = 1'b0;
      31'b0000000000000000000000000001000: n11902_o = 1'b0;
      31'b0000000000000000000000000000100: n11902_o = 1'b0;
      31'b0000000000000000000000000000010: n11902_o = 1'b0;
      31'b0000000000000000000000000000001: n11902_o = 1'b0;
      default: n11902_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11903_o = n10737_o;
      31'b0100000000000000000000000000000: n11903_o = n10737_o;
      31'b0010000000000000000000000000000: n11903_o = n10737_o;
      31'b0001000000000000000000000000000: n11903_o = n10737_o;
      31'b0000100000000000000000000000000: n11903_o = n10737_o;
      31'b0000010000000000000000000000000: n11903_o = n10737_o;
      31'b0000001000000000000000000000000: n11903_o = n11732_o;
      31'b0000000100000000000000000000000: n11903_o = n10737_o;
      31'b0000000010000000000000000000000: n11903_o = n10737_o;
      31'b0000000001000000000000000000000: n11903_o = n10737_o;
      31'b0000000000100000000000000000000: n11903_o = n11547_o;
      31'b0000000000010000000000000000000: n11903_o = n10737_o;
      31'b0000000000001000000000000000000: n11903_o = n10737_o;
      31'b0000000000000100000000000000000: n11903_o = n10737_o;
      31'b0000000000000010000000000000000: n11903_o = n10737_o;
      31'b0000000000000001000000000000000: n11903_o = n10737_o;
      31'b0000000000000000100000000000000: n11903_o = n10737_o;
      31'b0000000000000000010000000000000: n11903_o = n10737_o;
      31'b0000000000000000001000000000000: n11903_o = n10737_o;
      31'b0000000000000000000100000000000: n11903_o = n10737_o;
      31'b0000000000000000000010000000000: n11903_o = n10737_o;
      31'b0000000000000000000001000000000: n11903_o = n10737_o;
      31'b0000000000000000000000100000000: n11903_o = n10737_o;
      31'b0000000000000000000000010000000: n11903_o = n10737_o;
      31'b0000000000000000000000001000000: n11903_o = n10737_o;
      31'b0000000000000000000000000100000: n11903_o = n10737_o;
      31'b0000000000000000000000000010000: n11903_o = n10737_o;
      31'b0000000000000000000000000001000: n11903_o = n10737_o;
      31'b0000000000000000000000000000100: n11903_o = n10737_o;
      31'b0000000000000000000000000000010: n11903_o = n10737_o;
      31'b0000000000000000000000000000001: n11903_o = n10737_o;
      default: n11903_o = n10737_o;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11906_o = n11060_o;
      31'b0100000000000000000000000000000: n11906_o = n11060_o;
      31'b0010000000000000000000000000000: n11906_o = n11060_o;
      31'b0001000000000000000000000000000: n11906_o = n11060_o;
      31'b0000100000000000000000000000000: n11906_o = n11060_o;
      31'b0000010000000000000000000000000: n11906_o = n11060_o;
      31'b0000001000000000000000000000000: n11906_o = n11060_o;
      31'b0000000100000000000000000000000: n11906_o = n11060_o;
      31'b0000000010000000000000000000000: n11906_o = n11060_o;
      31'b0000000001000000000000000000000: n11906_o = n11060_o;
      31'b0000000000100000000000000000000: n11906_o = n11060_o;
      31'b0000000000010000000000000000000: n11906_o = n11060_o;
      31'b0000000000001000000000000000000: n11906_o = n11060_o;
      31'b0000000000000100000000000000000: n11906_o = n11060_o;
      31'b0000000000000010000000000000000: n11906_o = n11060_o;
      31'b0000000000000001000000000000000: n11906_o = n11060_o;
      31'b0000000000000000100000000000000: n11906_o = n11060_o;
      31'b0000000000000000010000000000000: n11906_o = n11060_o;
      31'b0000000000000000001000000000000: n11906_o = n11060_o;
      31'b0000000000000000000100000000000: n11906_o = n11060_o;
      31'b0000000000000000000010000000000: n11906_o = n11060_o;
      31'b0000000000000000000001000000000: n11906_o = n11060_o;
      31'b0000000000000000000000100000000: n11906_o = n11060_o;
      31'b0000000000000000000000010000000: n11906_o = n11060_o;
      31'b0000000000000000000000001000000: n11906_o = n11192_o;
      31'b0000000000000000000000000100000: n11906_o = n11060_o;
      31'b0000000000000000000000000010000: n11906_o = n11060_o;
      31'b0000000000000000000000000001000: n11906_o = n11060_o;
      31'b0000000000000000000000000000100: n11906_o = n11060_o;
      31'b0000000000000000000000000000010: n11906_o = n11104_o;
      31'b0000000000000000000000000000001: n11906_o = n11060_o;
      default: n11906_o = n11060_o;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11909_o = 1'b0;
      31'b0100000000000000000000000000000: n11909_o = 1'b0;
      31'b0010000000000000000000000000000: n11909_o = 1'b0;
      31'b0001000000000000000000000000000: n11909_o = 1'b0;
      31'b0000100000000000000000000000000: n11909_o = 1'b0;
      31'b0000010000000000000000000000000: n11909_o = 1'b0;
      31'b0000001000000000000000000000000: n11909_o = n11734_o;
      31'b0000000100000000000000000000000: n11909_o = 1'b0;
      31'b0000000010000000000000000000000: n11909_o = 1'b0;
      31'b0000000001000000000000000000000: n11909_o = 1'b0;
      31'b0000000000100000000000000000000: n11909_o = n11549_o;
      31'b0000000000010000000000000000000: n11909_o = 1'b0;
      31'b0000000000001000000000000000000: n11909_o = 1'b0;
      31'b0000000000000100000000000000000: n11909_o = 1'b0;
      31'b0000000000000010000000000000000: n11909_o = 1'b0;
      31'b0000000000000001000000000000000: n11909_o = 1'b0;
      31'b0000000000000000100000000000000: n11909_o = 1'b0;
      31'b0000000000000000010000000000000: n11909_o = 1'b0;
      31'b0000000000000000001000000000000: n11909_o = 1'b0;
      31'b0000000000000000000100000000000: n11909_o = 1'b0;
      31'b0000000000000000000010000000000: n11909_o = 1'b0;
      31'b0000000000000000000001000000000: n11909_o = 1'b0;
      31'b0000000000000000000000100000000: n11909_o = 1'b0;
      31'b0000000000000000000000010000000: n11909_o = 1'b0;
      31'b0000000000000000000000001000000: n11909_o = 1'b0;
      31'b0000000000000000000000000100000: n11909_o = 1'b0;
      31'b0000000000000000000000000010000: n11909_o = 1'b0;
      31'b0000000000000000000000000001000: n11909_o = 1'b0;
      31'b0000000000000000000000000000100: n11909_o = n11117_o;
      31'b0000000000000000000000000000010: n11909_o = n11107_o;
      31'b0000000000000000000000000000001: n11909_o = 1'b1;
      default: n11909_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11913_o = 1'b0;
      31'b0100000000000000000000000000000: n11913_o = 1'b0;
      31'b0010000000000000000000000000000: n11913_o = 1'b0;
      31'b0001000000000000000000000000000: n11913_o = 1'b0;
      31'b0000100000000000000000000000000: n11913_o = 1'b0;
      31'b0000010000000000000000000000000: n11913_o = 1'b0;
      31'b0000001000000000000000000000000: n11913_o = 1'b0;
      31'b0000000100000000000000000000000: n11913_o = 1'b0;
      31'b0000000010000000000000000000000: n11913_o = 1'b0;
      31'b0000000001000000000000000000000: n11913_o = 1'b0;
      31'b0000000000100000000000000000000: n11913_o = 1'b0;
      31'b0000000000010000000000000000000: n11913_o = 1'b0;
      31'b0000000000001000000000000000000: n11913_o = 1'b0;
      31'b0000000000000100000000000000000: n11913_o = 1'b0;
      31'b0000000000000010000000000000000: n11913_o = 1'b0;
      31'b0000000000000001000000000000000: n11913_o = 1'b0;
      31'b0000000000000000100000000000000: n11913_o = 1'b0;
      31'b0000000000000000010000000000000: n11913_o = 1'b1;
      31'b0000000000000000001000000000000: n11913_o = n11304_o;
      31'b0000000000000000000100000000000: n11913_o = 1'b1;
      31'b0000000000000000000010000000000: n11913_o = 1'b0;
      31'b0000000000000000000001000000000: n11913_o = 1'b0;
      31'b0000000000000000000000100000000: n11913_o = 1'b0;
      31'b0000000000000000000000010000000: n11913_o = 1'b0;
      31'b0000000000000000000000001000000: n11913_o = 1'b0;
      31'b0000000000000000000000000100000: n11913_o = 1'b0;
      31'b0000000000000000000000000010000: n11913_o = 1'b0;
      31'b0000000000000000000000000001000: n11913_o = 1'b0;
      31'b0000000000000000000000000000100: n11913_o = 1'b0;
      31'b0000000000000000000000000000010: n11913_o = 1'b0;
      31'b0000000000000000000000000000001: n11913_o = 1'b0;
      default: n11913_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11916_o = 1'b0;
      31'b0100000000000000000000000000000: n11916_o = 1'b0;
      31'b0010000000000000000000000000000: n11916_o = 1'b0;
      31'b0001000000000000000000000000000: n11916_o = 1'b0;
      31'b0000100000000000000000000000000: n11916_o = 1'b0;
      31'b0000010000000000000000000000000: n11916_o = 1'b0;
      31'b0000001000000000000000000000000: n11916_o = 1'b0;
      31'b0000000100000000000000000000000: n11916_o = 1'b0;
      31'b0000000010000000000000000000000: n11916_o = 1'b0;
      31'b0000000001000000000000000000000: n11916_o = 1'b0;
      31'b0000000000100000000000000000000: n11916_o = 1'b0;
      31'b0000000000010000000000000000000: n11916_o = 1'b0;
      31'b0000000000001000000000000000000: n11916_o = 1'b0;
      31'b0000000000000100000000000000000: n11916_o = 1'b0;
      31'b0000000000000010000000000000000: n11916_o = 1'b0;
      31'b0000000000000001000000000000000: n11916_o = 1'b0;
      31'b0000000000000000100000000000000: n11916_o = 1'b0;
      31'b0000000000000000010000000000000: n11916_o = 1'b0;
      31'b0000000000000000001000000000000: n11916_o = n11306_o;
      31'b0000000000000000000100000000000: n11916_o = 1'b1;
      31'b0000000000000000000010000000000: n11916_o = 1'b0;
      31'b0000000000000000000001000000000: n11916_o = 1'b0;
      31'b0000000000000000000000100000000: n11916_o = 1'b0;
      31'b0000000000000000000000010000000: n11916_o = 1'b0;
      31'b0000000000000000000000001000000: n11916_o = 1'b0;
      31'b0000000000000000000000000100000: n11916_o = 1'b0;
      31'b0000000000000000000000000010000: n11916_o = 1'b0;
      31'b0000000000000000000000000001000: n11916_o = 1'b0;
      31'b0000000000000000000000000000100: n11916_o = 1'b0;
      31'b0000000000000000000000000000010: n11916_o = 1'b0;
      31'b0000000000000000000000000000001: n11916_o = 1'b0;
      default: n11916_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11920_o = 1'b0;
      31'b0100000000000000000000000000000: n11920_o = 1'b0;
      31'b0010000000000000000000000000000: n11920_o = 1'b0;
      31'b0001000000000000000000000000000: n11920_o = 1'b0;
      31'b0000100000000000000000000000000: n11920_o = 1'b0;
      31'b0000010000000000000000000000000: n11920_o = 1'b0;
      31'b0000001000000000000000000000000: n11920_o = 1'b0;
      31'b0000000100000000000000000000000: n11920_o = 1'b0;
      31'b0000000010000000000000000000000: n11920_o = 1'b0;
      31'b0000000001000000000000000000000: n11920_o = 1'b0;
      31'b0000000000100000000000000000000: n11920_o = 1'b0;
      31'b0000000000010000000000000000000: n11920_o = 1'b0;
      31'b0000000000001000000000000000000: n11920_o = 1'b0;
      31'b0000000000000100000000000000000: n11920_o = 1'b0;
      31'b0000000000000010000000000000000: n11920_o = 1'b0;
      31'b0000000000000001000000000000000: n11920_o = 1'b0;
      31'b0000000000000000100000000000000: n11920_o = 1'b0;
      31'b0000000000000000010000000000000: n11920_o = 1'b1;
      31'b0000000000000000001000000000000: n11920_o = n11287_o;
      31'b0000000000000000000100000000000: n11920_o = 1'b1;
      31'b0000000000000000000010000000000: n11920_o = 1'b0;
      31'b0000000000000000000001000000000: n11920_o = 1'b0;
      31'b0000000000000000000000100000000: n11920_o = 1'b0;
      31'b0000000000000000000000010000000: n11920_o = 1'b0;
      31'b0000000000000000000000001000000: n11920_o = 1'b0;
      31'b0000000000000000000000000100000: n11920_o = 1'b0;
      31'b0000000000000000000000000010000: n11920_o = 1'b0;
      31'b0000000000000000000000000001000: n11920_o = 1'b0;
      31'b0000000000000000000000000000100: n11920_o = 1'b0;
      31'b0000000000000000000000000000010: n11920_o = 1'b0;
      31'b0000000000000000000000000000001: n11920_o = 1'b0;
      default: n11920_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11923_o = 1'b0;
      31'b0100000000000000000000000000000: n11923_o = 1'b0;
      31'b0010000000000000000000000000000: n11923_o = 1'b0;
      31'b0001000000000000000000000000000: n11923_o = 1'b0;
      31'b0000100000000000000000000000000: n11923_o = 1'b0;
      31'b0000010000000000000000000000000: n11923_o = 1'b0;
      31'b0000001000000000000000000000000: n11923_o = 1'b0;
      31'b0000000100000000000000000000000: n11923_o = 1'b0;
      31'b0000000010000000000000000000000: n11923_o = 1'b0;
      31'b0000000001000000000000000000000: n11923_o = 1'b0;
      31'b0000000000100000000000000000000: n11923_o = 1'b0;
      31'b0000000000010000000000000000000: n11923_o = 1'b0;
      31'b0000000000001000000000000000000: n11923_o = 1'b0;
      31'b0000000000000100000000000000000: n11923_o = 1'b0;
      31'b0000000000000010000000000000000: n11923_o = 1'b0;
      31'b0000000000000001000000000000000: n11923_o = 1'b0;
      31'b0000000000000000100000000000000: n11923_o = 1'b0;
      31'b0000000000000000010000000000000: n11923_o = 1'b1;
      31'b0000000000000000001000000000000: n11923_o = n11288_o;
      31'b0000000000000000000100000000000: n11923_o = n11224_o;
      31'b0000000000000000000010000000000: n11923_o = 1'b0;
      31'b0000000000000000000001000000000: n11923_o = 1'b0;
      31'b0000000000000000000000100000000: n11923_o = 1'b0;
      31'b0000000000000000000000010000000: n11923_o = 1'b0;
      31'b0000000000000000000000001000000: n11923_o = 1'b0;
      31'b0000000000000000000000000100000: n11923_o = 1'b0;
      31'b0000000000000000000000000010000: n11923_o = 1'b0;
      31'b0000000000000000000000000001000: n11923_o = 1'b0;
      31'b0000000000000000000000000000100: n11923_o = 1'b0;
      31'b0000000000000000000000000000010: n11923_o = 1'b0;
      31'b0000000000000000000000000000001: n11923_o = 1'b0;
      default: n11923_o = 1'b0;
    endcase
  /* execute1.vhdl:916:13  */
  always @*
    case (n11798_o)
      31'b1000000000000000000000000000000: n11927_o = n10832_o;
      31'b0100000000000000000000000000000: n11927_o = n10832_o;
      31'b0010000000000000000000000000000: n11927_o = n10832_o;
      31'b0001000000000000000000000000000: n11927_o = n10832_o;
      31'b0000100000000000000000000000000: n11927_o = n10832_o;
      31'b0000010000000000000000000000000: n11927_o = n10832_o;
      31'b0000001000000000000000000000000: n11927_o = n10832_o;
      31'b0000000100000000000000000000000: n11927_o = n10832_o;
      31'b0000000010000000000000000000000: n11927_o = n10832_o;
      31'b0000000001000000000000000000000: n11927_o = n10832_o;
      31'b0000000000100000000000000000000: n11927_o = n10832_o;
      31'b0000000000010000000000000000000: n11927_o = n10832_o;
      31'b0000000000001000000000000000000: n11927_o = n10832_o;
      31'b0000000000000100000000000000000: n11927_o = n10832_o;
      31'b0000000000000010000000000000000: n11927_o = n10832_o;
      31'b0000000000000001000000000000000: n11927_o = n10832_o;
      31'b0000000000000000100000000000000: n11927_o = n10832_o;
      31'b0000000000000000010000000000000: n11927_o = 1'b0;
      31'b0000000000000000001000000000000: n11927_o = n11301_o;
      31'b0000000000000000000100000000000: n11927_o = n11227_o;
      31'b0000000000000000000010000000000: n11927_o = n10832_o;
      31'b0000000000000000000001000000000: n11927_o = n10832_o;
      31'b0000000000000000000000100000000: n11927_o = n10832_o;
      31'b0000000000000000000000010000000: n11927_o = n10832_o;
      31'b0000000000000000000000001000000: n11927_o = n10832_o;
      31'b0000000000000000000000000100000: n11927_o = n10832_o;
      31'b0000000000000000000000000010000: n11927_o = n10832_o;
      31'b0000000000000000000000000001000: n11927_o = n10832_o;
      31'b0000000000000000000000000000100: n11927_o = n10832_o;
      31'b0000000000000000000000000000010: n11927_o = n10832_o;
      31'b0000000000000000000000000000001: n11927_o = n10832_o;
      default: n11927_o = n10832_o;
    endcase
  /* execute1.vhdl:1193:43  */
  assign n11928_o = n9139_o[73:10];
  assign n11929_o = ctrl[255:192];
  /* execute1.vhdl:1191:13  */
  assign n11930_o = n11941_o ? n11928_o : n11929_o;
  /* execute1.vhdl:1195:17  */
  assign n11932_o = n11920_o ? b_in : 64'b0000000000000000000000000000000000000000000000000000000000000100;
  assign n11933_o = n11886_o[2];
  /* execute1.vhdl:1195:17  */
  assign n11934_o = n11920_o ? n11923_o : n11933_o;
  /* execute1.vhdl:1201:41  */
  assign n11935_o = n9139_o[383];
  /* execute1.vhdl:1201:33  */
  assign n11936_o = n11920_o != n11935_o;
  /* execute1.vhdl:1191:13  */
  assign n11938_o = n11943_o ? 1'b1 : n11871_o;
  /* execute1.vhdl:1191:13  */
  assign n11939_o = n11947_o ? n11916_o : 1'b0;
  /* execute1.vhdl:1191:13  */
  assign n11941_o = n11913_o & n11920_o;
  assign n11942_o = {n11934_o, n11920_o, n11916_o, n11932_o};
  /* execute1.vhdl:1191:13  */
  assign n11943_o = n11913_o & n11936_o;
  assign n11944_o = n11886_o[2:0];
  assign n11945_o = {n11944_o, n11881_o};
  /* execute1.vhdl:1191:13  */
  assign n11946_o = n11913_o ? n11942_o : n11945_o;
  /* execute1.vhdl:1191:13  */
  assign n11947_o = n11913_o & n11936_o;
  assign n11948_o = n11886_o[3];
  /* execute1.vhdl:1209:44  */
  assign n11949_o = ~n11060_o;
  /* execute1.vhdl:1209:30  */
  assign n11950_o = valid_in & n11949_o;
  /* execute1.vhdl:1209:50  */
  assign n11952_o = n11950_o & 1'b1;
  /* execute1.vhdl:1211:21  */
  assign n11953_o = n9139_o[2:1];
  /* execute1.vhdl:1211:26  */
  assign n11955_o = n11953_o == 2'b10;
  /* execute1.vhdl:1213:24  */
  assign n11957_o = n9139_o[2:1];
  /* execute1.vhdl:1213:29  */
  assign n11959_o = n11957_o == 2'b00;
  /* execute1.vhdl:1215:36  */
  assign n11960_o = n9139_o[2:1];
  /* execute1.vhdl:1215:41  */
  assign n11962_o = n11960_o == 2'b11;
  /* execute1.vhdl:1215:27  */
  assign n11964_o = 1'b1 & n11962_o;
  /* execute1.vhdl:1215:13  */
  assign n11967_o = n11964_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:1213:13  */
  assign n11970_o = n11959_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:1213:13  */
  assign n11972_o = n11959_o ? 1'b0 : n11967_o;
  /* execute1.vhdl:1211:13  */
  assign n11974_o = n11955_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:1211:13  */
  assign n11976_o = n11955_o ? 1'b0 : n11970_o;
  /* execute1.vhdl:1211:13  */
  assign n11978_o = n11955_o ? 1'b0 : n11972_o;
  /* execute1.vhdl:1219:21  */
  assign n11979_o = n9139_o[9:4];
  /* execute1.vhdl:1219:31  */
  assign n11981_o = n11979_o == 6'b111101;
  /* execute1.vhdl:1209:9  */
  assign n11983_o = n11988_o ? 1'b0 : n10832_o;
  /* execute1.vhdl:1209:9  */
  assign n11985_o = n11952_o ? n11974_o : 1'b0;
  /* execute1.vhdl:1209:9  */
  assign n11987_o = n11952_o ? n11976_o : 1'b0;
  /* execute1.vhdl:1209:9  */
  assign n11988_o = n11952_o & n11981_o;
  /* execute1.vhdl:1209:9  */
  assign n11990_o = n11952_o ? n11978_o : 1'b0;
  /* execute1.vhdl:913:9  */
  assign n11992_o = n11094_o ? n11801_o : 1'b0;
  assign n11994_o = {n11930_o, n11846_o, n11843_o, n11840_o, n11836_o, n11833_o, n11830_o, n11827_o, n11825_o, n11822_o, n11819_o, n11815_o, n11812_o, n11808_o, n11805_o, n11802_o};
  assign n11995_o = {n10753_o, n10752_o};
  /* execute1.vhdl:913:9  */
  assign n11998_o = n11094_o ? n11848_o : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* execute1.vhdl:913:9  */
  assign n12000_o = n11094_o ? n11849_o : 1'b0;
  /* execute1.vhdl:913:9  */
  assign n12001_o = n11094_o ? n11850_o : 1'b0;
  assign n12002_o = {n11852_o, n11851_o};
  assign n12003_o = {1'b0, 1'b0};
  /* execute1.vhdl:913:9  */
  assign n12004_o = n11094_o ? n12002_o : n12003_o;
  assign n12005_o = {n11893_o, n11889_o, n11948_o, n11946_o, n11877_o, n11874_o, n11938_o, n11868_o, n11865_o, n11862_o, n11859_o, n11855_o};
  assign n12006_o = {n11895_o, n11894_o};
  assign n12007_o = {n11899_o, n11898_o};
  assign n12008_o = {n11901_o, n11900_o};
  assign n12009_o = {n11903_o, n11939_o, n11902_o};
  assign n12010_o = {n10817_o, n11056_o, n11031_o, n11059_o, n11027_o, n11053_o, n11023_o, n11047_o, n11019_o, n11041_o, n11015_o, n10823_o, n10822_o, n10715_o, n10815_o, n11011_o, n10816_o, xerc_in, n10826_o, n10825_o, n10829_o, n10828_o, n10830_o};
  assign n12012_o = {1'b0, n11065_o};
  assign n12014_o = r[749];
  /* execute1.vhdl:913:9  */
  assign n12015_o = n11094_o ? n11897_o : n12014_o;
  assign n12016_o = {1'b0, n10837_o};
  assign n12018_o = {1'b0, 1'b0};
  assign n12020_o = {n10737_o, 1'b0, 1'b0};
  /* execute1.vhdl:913:9  */
  assign n12021_o = n11094_o ? n12009_o : n12020_o;
  assign n12022_o = r[750];
  /* execute1.vhdl:913:9  */
  assign n12026_o = n11094_o ? 1'b0 : n11985_o;
  /* execute1.vhdl:913:9  */
  assign n12029_o = n11094_o ? n11906_o : n11060_o;
  /* execute1.vhdl:913:9  */
  assign n12030_o = n11094_o ? n11909_o : n11987_o;
  /* execute1.vhdl:913:9  */
  assign n12047_o = n11094_o ? n11927_o : n11983_o;
  /* execute1.vhdl:913:9  */
  assign n12049_o = n11094_o ? 1'b0 : n11990_o;
  /* execute1.vhdl:1227:14  */
  assign n12052_o = r[761];
  /* execute1.vhdl:1230:17  */
  assign n12054_o = r[758];
  /* execute1.vhdl:1230:44  */
  assign n12055_o = r[760];
  /* execute1.vhdl:1230:39  */
  assign n12056_o = n12054_o | n12055_o;
  /* execute1.vhdl:1231:19  */
  assign n12057_o = r[758];
  /* execute1.vhdl:1231:59  */
  assign n12058_o = multiply_to_x[0];
  /* execute1.vhdl:1231:41  */
  assign n12059_o = n12057_o & n12058_o;
  /* execute1.vhdl:1232:19  */
  assign n12060_o = r[760];
  /* execute1.vhdl:1232:58  */
  assign n12061_o = divider_to_x[0];
  /* execute1.vhdl:1232:41  */
  assign n12062_o = n12060_o & n12061_o;
  /* execute1.vhdl:1231:72  */
  assign n12063_o = n12059_o | n12062_o;
  /* execute1.vhdl:1233:22  */
  assign n12064_o = r[758];
  /* execute1.vhdl:1236:46  */
  assign n12065_o = divider_to_x[65];
  /* execute1.vhdl:1233:17  */
  assign n12067_o = n12064_o ? 1'b0 : n12065_o;
  /* execute1.vhdl:1238:22  */
  assign n12068_o = r[758];
  /* execute1.vhdl:1238:56  */
  assign n12069_o = current[331];
  /* execute1.vhdl:1238:44  */
  assign n12070_o = n12068_o & n12069_o;
  /* execute1.vhdl:1246:32  */
  assign n12073_o = current[331];
  assign n12075_o = n12005_o[124];
  assign n12076_o = n12010_o[124];
  /* execute1.vhdl:913:9  */
  assign n12077_o = n11094_o ? n12075_o : n12076_o;
  /* execute1.vhdl:1249:25  */
  assign n12078_o = n12067_o ? 1'b1 : n12077_o;
  assign n12079_o = {n12078_o, n12067_o, n12067_o};
  assign n12080_o = n12005_o[124:122];
  assign n12081_o = n12010_o[124:122];
  /* execute1.vhdl:913:9  */
  assign n12082_o = n11094_o ? n12080_o : n12081_o;
  /* execute1.vhdl:1246:21  */
  assign n12083_o = n12073_o ? n12079_o : n12082_o;
  assign n12085_o = n12005_o[0];
  assign n12086_o = n12010_o[0];
  /* execute1.vhdl:913:9  */
  assign n12087_o = n11094_o ? n12085_o : n12086_o;
  /* execute1.vhdl:1238:17  */
  assign n12088_o = n12070_o ? n12087_o : 1'b1;
  assign n12089_o = n12005_o[124:122];
  assign n12090_o = n12010_o[124:122];
  /* execute1.vhdl:913:9  */
  assign n12091_o = n11094_o ? n12089_o : n12090_o;
  /* execute1.vhdl:1238:17  */
  assign n12092_o = n12070_o ? n12091_o : n12083_o;
  assign n12093_o = n12006_o[0];
  assign n12094_o = n12012_o[0];
  /* execute1.vhdl:913:9  */
  assign n12095_o = n11094_o ? n12093_o : n12094_o;
  /* execute1.vhdl:1238:17  */
  assign n12096_o = n12070_o ? 1'b1 : n12095_o;
  /* execute1.vhdl:1231:13  */
  assign n12097_o = n12114_o ? 1'b1 : 1'b0;
  /* execute1.vhdl:1257:40  */
  assign n12099_o = r[758];
  /* execute1.vhdl:1258:40  */
  assign n12100_o = r[760];
  assign n12101_o = n12005_o[0];
  assign n12102_o = n12010_o[0];
  /* execute1.vhdl:913:9  */
  assign n12103_o = n11094_o ? n12101_o : n12102_o;
  /* execute1.vhdl:1231:13  */
  assign n12104_o = n12063_o ? n12088_o : n12103_o;
  assign n12105_o = n12005_o[124:122];
  assign n12106_o = n12010_o[124:122];
  /* execute1.vhdl:913:9  */
  assign n12107_o = n11094_o ? n12105_o : n12106_o;
  /* execute1.vhdl:1231:13  */
  assign n12108_o = n12063_o ? n12092_o : n12107_o;
  /* execute1.vhdl:1231:13  */
  assign n12109_o = n12063_o ? n12096_o : 1'b1;
  assign n12110_o = n12007_o[1];
  assign n12111_o = n12016_o[1];
  /* execute1.vhdl:913:9  */
  assign n12112_o = n11094_o ? n12110_o : n12111_o;
  /* execute1.vhdl:1231:13  */
  assign n12113_o = n12063_o ? n12112_o : n12099_o;
  /* execute1.vhdl:1231:13  */
  assign n12114_o = n12063_o & n12070_o;
  assign n12115_o = n12008_o[0];
  assign n12116_o = n12018_o[0];
  /* execute1.vhdl:913:9  */
  assign n12117_o = n11094_o ? n12115_o : n12116_o;
  /* execute1.vhdl:1231:13  */
  assign n12118_o = n12063_o ? n12117_o : n12100_o;
  /* execute1.vhdl:1260:17  */
  assign n12120_o = r[759];
  /* execute1.vhdl:1262:42  */
  assign n12121_o = multiply_to_x[129];
  /* execute1.vhdl:1263:44  */
  assign n12122_o = multiply_to_x[129];
  /* execute1.vhdl:1264:30  */
  assign n12123_o = multiply_to_x[129];
  assign n12125_o = n12005_o[124];
  assign n12126_o = n12010_o[124];
  /* execute1.vhdl:913:9  */
  assign n12127_o = n11094_o ? n12125_o : n12126_o;
  /* execute1.vhdl:1264:13  */
  assign n12128_o = n12123_o ? 1'b1 : n12127_o;
  assign n12130_o = {n12128_o, n12122_o, n12121_o};
  assign n12131_o = n12005_o[0];
  assign n12132_o = n12010_o[0];
  /* execute1.vhdl:913:9  */
  assign n12133_o = n11094_o ? n12131_o : n12132_o;
  /* execute1.vhdl:1260:9  */
  assign n12134_o = n12120_o ? 1'b1 : n12133_o;
  assign n12135_o = n12005_o[124:122];
  assign n12136_o = n12010_o[124:122];
  /* execute1.vhdl:913:9  */
  assign n12137_o = n11094_o ? n12135_o : n12136_o;
  /* execute1.vhdl:1260:9  */
  assign n12138_o = n12120_o ? n12130_o : n12137_o;
  /* execute1.vhdl:1260:9  */
  assign n12141_o = n12120_o ? 1'b1 : 1'b0;
  assign n12142_o = {n12118_o, n12097_o, n12113_o};
  /* execute1.vhdl:1230:9  */
  assign n12143_o = n12056_o ? n12104_o : n12134_o;
  /* execute1.vhdl:1230:9  */
  assign n12144_o = n12056_o ? n12108_o : n12138_o;
  assign n12145_o = n12006_o[0];
  assign n12146_o = n12012_o[0];
  /* execute1.vhdl:913:9  */
  assign n12147_o = n11094_o ? n12145_o : n12146_o;
  /* execute1.vhdl:1230:9  */
  assign n12148_o = n12056_o ? n12109_o : n12147_o;
  assign n12149_o = n12007_o[1];
  assign n12150_o = n12016_o[1];
  /* execute1.vhdl:913:9  */
  assign n12151_o = n11094_o ? n12149_o : n12150_o;
  assign n12152_o = n12008_o[0];
  assign n12153_o = n12018_o[0];
  /* execute1.vhdl:913:9  */
  assign n12154_o = n11094_o ? n12152_o : n12153_o;
  assign n12155_o = {n12154_o, 1'b0, n12151_o};
  /* execute1.vhdl:1230:9  */
  assign n12156_o = n12056_o ? n12142_o : n12155_o;
  /* execute1.vhdl:1230:9  */
  assign n12159_o = n12056_o ? 1'b0 : n12141_o;
  /* execute1.vhdl:1227:9  */
  assign n12160_o = n12052_o ? 1'b1 : n12143_o;
  assign n12161_o = n12005_o[124:122];
  assign n12162_o = n12010_o[124:122];
  /* execute1.vhdl:913:9  */
  assign n12163_o = n11094_o ? n12161_o : n12162_o;
  /* execute1.vhdl:1227:9  */
  assign n12164_o = n12052_o ? n12163_o : n12144_o;
  assign n12165_o = n12006_o[0];
  assign n12166_o = n12012_o[0];
  /* execute1.vhdl:913:9  */
  assign n12167_o = n11094_o ? n12165_o : n12166_o;
  /* execute1.vhdl:1227:9  */
  assign n12168_o = n12052_o ? n12167_o : n12148_o;
  assign n12169_o = n12007_o[1];
  assign n12170_o = n12016_o[1];
  /* execute1.vhdl:913:9  */
  assign n12171_o = n11094_o ? n12169_o : n12170_o;
  assign n12172_o = n12008_o[0];
  assign n12173_o = n12018_o[0];
  /* execute1.vhdl:913:9  */
  assign n12174_o = n11094_o ? n12172_o : n12173_o;
  assign n12175_o = {n12174_o, 1'b0, n12171_o};
  /* execute1.vhdl:1227:9  */
  assign n12176_o = n12052_o ? n12175_o : n12156_o;
  assign n12183_o = n12005_o[121:1];
  assign n12184_o = n12010_o[121:1];
  /* execute1.vhdl:913:9  */
  assign n12185_o = n11094_o ? n12183_o : n12184_o;
  assign n12186_o = n12006_o[1];
  assign n12187_o = n12012_o[1];
  /* execute1.vhdl:913:9  */
  assign n12188_o = n11094_o ? n12186_o : n12187_o;
  assign n12189_o = n12007_o[0];
  assign n12190_o = n12016_o[0];
  /* execute1.vhdl:913:9  */
  assign n12191_o = n11094_o ? n12189_o : n12190_o;
  assign n12192_o = n12008_o[1];
  assign n12193_o = n12018_o[1];
  /* execute1.vhdl:913:9  */
  assign n12194_o = n11094_o ? n12192_o : n12193_o;
  /* execute1.vhdl:1227:9  */
  assign n12197_o = n12052_o ? 1'b0 : n12159_o;
  assign n12201_o = n12005_o[137:126];
  assign n12202_o = n12010_o[137:126];
  /* execute1.vhdl:913:9  */
  assign n12203_o = n11094_o ? n12201_o : n12202_o;
  /* execute1.vhdl:1270:9  */
  assign n12204_o = n12030_o ? 12'b011100000000 : n12203_o;
  assign n12205_o = n12005_o[277];
  assign n12206_o = n12010_o[277];
  /* execute1.vhdl:913:9  */
  assign n12207_o = n11094_o ? n12205_o : n12206_o;
  /* execute1.vhdl:1270:9  */
  assign n12208_o = n12030_o ? 1'b1 : n12207_o;
  assign n12215_o = n12005_o[353:278];
  assign n12216_o = n12010_o[353:278];
  /* execute1.vhdl:913:9  */
  assign n12217_o = n11094_o ? n12215_o : n12216_o;
  assign n12218_o = n12005_o[276:138];
  assign n12219_o = n12010_o[276:138];
  /* execute1.vhdl:913:9  */
  assign n12220_o = n11094_o ? n12218_o : n12219_o;
  /* execute1.vhdl:1270:9  */
  assign n12222_o = n12030_o ? 1'b1 : n12029_o;
  /* execute1.vhdl:1279:50  */
  assign n12223_o = n9140_o[1];
  /* execute1.vhdl:1279:70  */
  assign n12224_o = n9140_o[2];
  /* execute1.vhdl:1279:62  */
  assign n12225_o = n12223_o | n12224_o;
  /* execute1.vhdl:1279:40  */
  assign n12226_o = ~n12225_o;
  /* execute1.vhdl:1279:36  */
  assign n12227_o = n12222_o & n12226_o;
  assign n12228_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12022_o, n12015_o, n11071_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12185_o, n12160_o};
  /* execute1.vhdl:1280:14  */
  assign n12229_o = n12228_o[353:0];
  /* execute1.vhdl:1280:16  */
  assign n12230_o = n12229_o[125];
  /* execute1.vhdl:1280:9  */
  assign n12232_o = n12230_o ? 1'b0 : n11071_o;
  /* execute1.vhdl:1284:9  */
  assign n12234_o = n12047_o ? 1'b1 : n12022_o;
  assign n12250_o = {1'b0, 1'b1};
  assign n12251_o = {1'b0, 1'b0};
  assign n12252_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n12253_o = {1'b0, 1'b0, 1'b0};
  assign n12254_o = n11994_o[65:64];
  assign n12255_o = n11995_o[65:64];
  /* execute1.vhdl:913:9  */
  assign n12256_o = n11094_o ? n12254_o : n12255_o;
  /* execute1.vhdl:1288:9  */
  assign n12257_o = interrupt_in ? n12250_o : n12256_o;
  assign n12258_o = n11994_o[69:68];
  assign n12259_o = n11995_o[69:68];
  /* execute1.vhdl:913:9  */
  assign n12260_o = n11094_o ? n12258_o : n12259_o;
  /* execute1.vhdl:1288:9  */
  assign n12261_o = interrupt_in ? n12251_o : n12260_o;
  assign n12262_o = n11994_o[75:72];
  assign n12263_o = n11995_o[75:72];
  /* execute1.vhdl:913:9  */
  assign n12264_o = n11094_o ? n12262_o : n12263_o;
  /* execute1.vhdl:1288:9  */
  assign n12265_o = interrupt_in ? n12252_o : n12264_o;
  assign n12266_o = n11994_o[79:77];
  assign n12267_o = n11995_o[79:77];
  /* execute1.vhdl:913:9  */
  assign n12268_o = n11094_o ? n12266_o : n12267_o;
  /* execute1.vhdl:1288:9  */
  assign n12269_o = interrupt_in ? n12253_o : n12268_o;
  assign n12270_o = n11994_o[127];
  assign n12271_o = n11995_o[127];
  /* execute1.vhdl:913:9  */
  assign n12272_o = n11094_o ? n12270_o : n12271_o;
  /* execute1.vhdl:1288:9  */
  assign n12273_o = interrupt_in ? 1'b1 : n12272_o;
  assign n12277_o = n11994_o[63:0];
  assign n12278_o = n11995_o[63:0];
  /* execute1.vhdl:913:9  */
  assign n12279_o = n11094_o ? n12277_o : n12278_o;
  assign n12283_o = n11994_o[67:66];
  assign n12284_o = n11995_o[67:66];
  /* execute1.vhdl:913:9  */
  assign n12285_o = n11094_o ? n12283_o : n12284_o;
  assign n12289_o = n11994_o[71:70];
  assign n12290_o = n11995_o[71:70];
  /* execute1.vhdl:913:9  */
  assign n12291_o = n11094_o ? n12289_o : n12290_o;
  assign n12295_o = n11994_o[76];
  assign n12296_o = n11995_o[76];
  /* execute1.vhdl:913:9  */
  assign n12297_o = n11094_o ? n12295_o : n12296_o;
  assign n12298_o = n11994_o[191:128];
  assign n12299_o = n11995_o[191:128];
  /* execute1.vhdl:913:9  */
  assign n12300_o = n11094_o ? n12298_o : n12299_o;
  assign n12301_o = n11994_o[126:80];
  assign n12302_o = n11995_o[126:80];
  /* execute1.vhdl:913:9  */
  assign n12303_o = n11094_o ? n12301_o : n12302_o;
  assign n12304_o = {1'b0, 1'b0, 1'b0};
  assign n12305_o = {n12234_o, n12015_o, n12232_o};
  /* execute1.vhdl:1288:9  */
  assign n12306_o = interrupt_in ? n12304_o : n12305_o;
  /* execute1.vhdl:1306:25  */
  assign n12307_o = ~n12197_o;
  /* execute1.vhdl:1309:33  */
  assign n12308_o = r[353:0];
  /* execute1.vhdl:1309:35  */
  assign n12309_o = n12308_o[77:14];
  /* execute1.vhdl:1306:9  */
  assign n12310_o = n12307_o ? alu_result : n12309_o;
  assign n12311_o = n12005_o[121:78];
  assign n12312_o = n12010_o[121:78];
  /* execute1.vhdl:913:9  */
  assign n12313_o = n11094_o ? n12311_o : n12312_o;
  /* execute1.vhdl:1311:34  */
  assign n12317_o = current[83:77];
  assign n12318_o = n12005_o[6:1];
  assign n12319_o = n12010_o[6:1];
  /* execute1.vhdl:913:9  */
  assign n12320_o = n11094_o ? n12318_o : n12319_o;
  /* execute1.vhdl:1312:37  */
  assign n12321_o = current[84];
  assign n12322_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12313_o, n12310_o, n12317_o, n12320_o, n12160_o};
  /* execute1.vhdl:1312:60  */
  assign n12323_o = n12322_o[353:0];
  /* execute1.vhdl:1312:62  */
  assign n12324_o = n12323_o[0];
  /* execute1.vhdl:1312:54  */
  assign n12325_o = n12321_o & n12324_o;
  /* execute1.vhdl:1312:72  */
  assign n12326_o = ~n12222_o;
  /* execute1.vhdl:1312:68  */
  assign n12327_o = n12325_o & n12326_o;
  assign n12328_o = n12005_o[5:1];
  assign n12329_o = n12010_o[5:1];
  /* execute1.vhdl:913:9  */
  assign n12330_o = n11094_o ? n12328_o : n12329_o;
  /* execute1.vhdl:1313:27  */
  assign n12331_o = current[330];
  assign n12332_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12313_o, n12310_o, n12317_o, n12327_o, n12330_o, n12160_o};
  /* execute1.vhdl:1313:36  */
  assign n12333_o = n12332_o[353:0];
  /* execute1.vhdl:1313:38  */
  assign n12334_o = n12333_o[0];
  /* execute1.vhdl:1313:30  */
  assign n12335_o = n12331_o & n12334_o;
  /* execute1.vhdl:1313:48  */
  assign n12336_o = ~n12222_o;
  /* execute1.vhdl:1313:44  */
  assign n12337_o = n12335_o & n12336_o;
  assign n12338_o = n12005_o[5];
  assign n12339_o = n12010_o[5];
  /* execute1.vhdl:913:9  */
  assign n12340_o = n11094_o ? n12338_o : n12339_o;
  assign n12341_o = n12005_o[3:1];
  assign n12342_o = n12010_o[3:1];
  /* execute1.vhdl:913:9  */
  assign n12343_o = n11094_o ? n12341_o : n12342_o;
  assign n12344_o = n12005_o[121:119];
  assign n12345_o = n12010_o[121:119];
  /* execute1.vhdl:913:9  */
  assign n12346_o = n11094_o ? n12344_o : n12345_o;
  assign n12350_o = n12005_o[78];
  assign n12351_o = n12010_o[78];
  /* execute1.vhdl:913:9  */
  assign n12352_o = n11094_o ? n12350_o : n12351_o;
  /* execute1.vhdl:1316:40  */
  assign n12353_o = current[339];
  assign n12354_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12346_o, write_cr_data, write_cr_mask, n12352_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1316:56  */
  assign n12355_o = n12354_o[353:0];
  /* execute1.vhdl:1316:58  */
  assign n12356_o = n12355_o[0];
  /* execute1.vhdl:1316:50  */
  assign n12357_o = n12353_o & n12356_o;
  /* execute1.vhdl:1316:68  */
  assign n12358_o = ~n12222_o;
  /* execute1.vhdl:1316:64  */
  assign n12359_o = n12357_o & n12358_o;
  /* execute1.vhdl:1317:42  */
  assign n12360_o = current[340];
  assign n12361_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12346_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1317:59  */
  assign n12362_o = n12361_o[353:0];
  /* execute1.vhdl:1317:61  */
  assign n12363_o = n12362_o[0];
  /* execute1.vhdl:1317:53  */
  assign n12364_o = n12360_o & n12363_o;
  /* execute1.vhdl:1317:71  */
  assign n12365_o = ~n12222_o;
  /* execute1.vhdl:1317:67  */
  assign n12366_o = n12364_o & n12365_o;
  assign n12367_o = n12005_o[121:120];
  assign n12368_o = n12010_o[121:120];
  /* execute1.vhdl:913:9  */
  assign n12369_o = n11094_o ? n12367_o : n12368_o;
  /* execute1.vhdl:1319:42  */
  assign n12370_o = current[76:74];
  /* execute1.vhdl:1319:52  */
  assign n12371_o = n12370_o[2];
  /* execute1.vhdl:1319:70  */
  assign n12372_o = current[84];
  /* execute1.vhdl:1319:58  */
  assign n12373_o = n12371_o & n12372_o;
  assign n12374_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1319:93  */
  assign n12375_o = n12374_o[353:0];
  /* execute1.vhdl:1319:95  */
  assign n12376_o = n12375_o[0];
  /* execute1.vhdl:1319:87  */
  assign n12377_o = n12373_o & n12376_o;
  /* execute1.vhdl:1320:40  */
  assign n12378_o = current[76:74];
  /* execute1.vhdl:1320:50  */
  assign n12379_o = n12378_o[1:0];
  assign n12380_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1321:31  */
  assign n12381_o = n12380_o[353:0];
  /* execute1.vhdl:1321:33  */
  assign n12382_o = n12381_o[77:14];
  /* execute1.vhdl:1323:45  */
  assign n12383_o = current[76:74];
  /* execute1.vhdl:1323:55  */
  assign n12384_o = n12383_o[2];
  /* execute1.vhdl:1323:73  */
  assign n12385_o = current[339];
  /* execute1.vhdl:1323:61  */
  assign n12386_o = n12384_o & n12385_o;
  assign n12387_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1323:89  */
  assign n12388_o = n12387_o[353:0];
  /* execute1.vhdl:1323:91  */
  assign n12389_o = n12388_o[0];
  /* execute1.vhdl:1323:83  */
  assign n12390_o = n12386_o & n12389_o;
  /* execute1.vhdl:1324:43  */
  assign n12391_o = current[76:74];
  /* execute1.vhdl:1324:53  */
  assign n12392_o = n12391_o[1:0];
  assign n12393_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1326:33  */
  assign n12394_o = n12393_o[79];
  assign n12395_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1327:77  */
  assign n12396_o = n12395_o[90:87];
  /* execute1.vhdl:1329:65  */
  assign n12397_o = cr_in[3:0];
  /* execute1.vhdl:1326:13  */
  assign n12398_o = n12394_o ? n12396_o : n12397_o;
  assign n12399_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1326:33  */
  assign n12400_o = n12399_o[80];
  assign n12401_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1327:77  */
  assign n12402_o = n12401_o[94:91];
  /* execute1.vhdl:1329:65  */
  assign n12403_o = cr_in[7:4];
  /* execute1.vhdl:1326:13  */
  assign n12404_o = n12400_o ? n12402_o : n12403_o;
  assign n12405_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1326:33  */
  assign n12406_o = n12405_o[81];
  assign n12407_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1327:77  */
  assign n12408_o = n12407_o[98:95];
  /* execute1.vhdl:1329:65  */
  assign n12409_o = cr_in[11:8];
  /* execute1.vhdl:1326:13  */
  assign n12410_o = n12406_o ? n12408_o : n12409_o;
  assign n12411_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1326:33  */
  assign n12412_o = n12411_o[82];
  assign n12413_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1327:77  */
  assign n12414_o = n12413_o[102:99];
  /* execute1.vhdl:1329:65  */
  assign n12415_o = cr_in[15:12];
  /* execute1.vhdl:1326:13  */
  assign n12416_o = n12412_o ? n12414_o : n12415_o;
  assign n12417_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1326:33  */
  assign n12418_o = n12417_o[83];
  assign n12419_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1327:77  */
  assign n12420_o = n12419_o[106:103];
  /* execute1.vhdl:1329:65  */
  assign n12421_o = cr_in[19:16];
  /* execute1.vhdl:1326:13  */
  assign n12422_o = n12418_o ? n12420_o : n12421_o;
  assign n12423_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1326:33  */
  assign n12424_o = n12423_o[84];
  assign n12425_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1327:77  */
  assign n12426_o = n12425_o[110:107];
  /* execute1.vhdl:1329:65  */
  assign n12427_o = cr_in[23:20];
  /* execute1.vhdl:1326:13  */
  assign n12428_o = n12424_o ? n12426_o : n12427_o;
  assign n12429_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1326:33  */
  assign n12430_o = n12429_o[85];
  assign n12431_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1327:77  */
  assign n12432_o = n12431_o[114:111];
  /* execute1.vhdl:1329:65  */
  assign n12433_o = cr_in[27:24];
  /* execute1.vhdl:1326:13  */
  assign n12434_o = n12430_o ? n12432_o : n12433_o;
  assign n12435_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1326:33  */
  assign n12436_o = n12435_o[86];
  assign n12437_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  /* execute1.vhdl:1327:77  */
  assign n12438_o = n12437_o[118:115];
  /* execute1.vhdl:1329:65  */
  assign n12439_o = cr_in[31:28];
  /* execute1.vhdl:1326:13  */
  assign n12440_o = n12436_o ? n12438_o : n12439_o;
  /* execute1.vhdl:1334:23  */
  assign n12441_o = n9139_o[9:4];
  /* execute1.vhdl:1335:24  */
  assign n12443_o = n9139_o[73:10];
  /* execute1.vhdl:1336:30  */
  assign n12445_o = n9139_o[76:74];
  /* execute1.vhdl:1340:30  */
  assign n12451_o = n9139_o[83:77];
  /* execute1.vhdl:1341:27  */
  assign n12453_o = n9139_o[378:375];
  /* execute1.vhdl:1342:33  */
  assign n12455_o = n9139_o[379];
  /* execute1.vhdl:1342:59  */
  assign n12456_o = ctrl[128];
  /* execute1.vhdl:1342:46  */
  assign n12457_o = ~(n12455_o ^ n12456_o);
  assign n12459_o = n12027_o[309];
  /* execute1.vhdl:1343:32  */
  assign n12460_o = n9139_o[380];
  /* execute1.vhdl:1344:27  */
  assign n12462_o = n9139_o[381];
  /* execute1.vhdl:1346:28  */
  assign n12465_o = n9139_o[382];
  /* execute1.vhdl:1347:23  */
  assign n12467_o = n9139_o[330];
  /* execute1.vhdl:1348:25  */
  assign n12469_o = n9139_o[374:343];
  /* execute1.vhdl:1350:21  */
  assign n12470_o = n9139_o[374:369];
  /* execute1.vhdl:1350:36  */
  assign n12472_o = n12470_o == 6'b011111;
  /* execute1.vhdl:1350:60  */
  assign n12473_o = n9139_o[353:352];
  /* execute1.vhdl:1350:74  */
  assign n12475_o = n12473_o == 2'b11;
  /* execute1.vhdl:1350:47  */
  assign n12476_o = n12472_o & n12475_o;
  /* execute1.vhdl:1351:22  */
  assign n12477_o = n9139_o[348:344];
  /* execute1.vhdl:1351:35  */
  assign n12479_o = n12477_o == 5'b10101;
  /* execute1.vhdl:1350:81  */
  assign n12480_o = n12476_o & n12479_o;
  /* execute1.vhdl:1350:9  */
  assign n12482_o = n12480_o ? 1'b1 : n12459_o;
  /* execute1.vhdl:1354:33  */
  assign n12483_o = ctrl[132];
  /* execute1.vhdl:1355:37  */
  assign n12485_o = ctrl[142];
  /* execute1.vhdl:1355:25  */
  assign n12486_o = ~n12485_o;
  /* execute1.vhdl:1356:38  */
  assign n12488_o = ctrl[191];
  /* execute1.vhdl:1356:26  */
  assign n12489_o = ~n12488_o;
  /* execute1.vhdl:1357:29  */
  assign n12491_o = n9139_o[341];
  /* execute1.vhdl:1358:27  */
  assign n12493_o = n9139_o[390];
  /* execute1.vhdl:1359:27  */
  assign n12495_o = n9139_o[391];
  assign n12496_o = n12027_o[389:326];
  /* execute1.vhdl:1362:23  */
  assign n12497_o = n9139_o[9:4];
  /* execute1.vhdl:1363:24  */
  assign n12499_o = n9139_o[73:10];
  /* execute1.vhdl:1364:25  */
  assign n12501_o = n9139_o[374:343];
  /* execute1.vhdl:1365:25  */
  assign n12504_o = n9139_o[76:74];
  /* execute1.vhdl:1366:27  */
  assign n12505_o = n9139_o[341];
  /* execute1.vhdl:1367:31  */
  assign n12507_o = ctrl[139];
  /* execute1.vhdl:1367:51  */
  assign n12508_o = ctrl[136];
  /* execute1.vhdl:1367:41  */
  assign n12509_o = {n12507_o, n12508_o};
  /* execute1.vhdl:1371:24  */
  assign n12514_o = n9139_o[83:77];
  /* execute1.vhdl:1372:23  */
  assign n12516_o = n9139_o[330];
  /* execute1.vhdl:1373:27  */
  assign n12518_o = n9139_o[339];
  assign n12519_o = {n12021_o, n11032_o, n11086_o, n11081_o, n12194_o, n12176_o, n12191_o, n10836_o, n12306_o, n12188_o, n12168_o, n10834_o, n12217_o, n12208_o, n12220_o, n12204_o, n12227_o, n12164_o, n12369_o, n12366_o, write_cr_data, write_cr_mask, n12359_o, n12310_o, n12317_o, n12327_o, n12340_o, n12337_o, n12343_o, n12160_o};
  assign n12520_o = {n12496_o, n12495_o, n12493_o, n12491_o, n12489_o, n12486_o, n12483_o, n12467_o, n12465_o, xerc_in, n12462_o, n12460_o, n12457_o, n12482_o, n12453_o, n12451_o, c_in, b_in, a_in, n12445_o, n12469_o, n12443_o, n12441_o, n12026_o};
  /* execute1.vhdl:1381:36  */
  assign n12523_o = ctrl[191:128];
  /* execute1.vhdl:230:37  */
  assign n12529_o = n12523_o[63:31];
  /* execute1.vhdl:231:37  */
  assign n12532_o = n12523_o[26:22];
  assign n12533_o = n12530_o[30:27];
  /* execute1.vhdl:232:37  */
  assign n12535_o = n12523_o[15:0];
  assign n12536_o = n12530_o[21:16];
  assign n12537_o = {n12529_o, n12533_o, n12532_o, n12536_o, n12535_o};
  assign n12538_o = r[289:0];
  assign n12539_o = {n12518_o, n12516_o, n12514_o, c_in, b_in, a_in, n12509_o, n12505_o, n12501_o, n12504_o, n12499_o, n12497_o, n12049_o};
  /* execute1.vhdl:404:9  */
  always @(posedge clk)
    n12548_q <= n9370_o;
  /* execute1.vhdl:404:9  */
  always @(posedge clk)
    n12549_q <= n9378_o;
  initial
    n12549_q = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* execute1.vhdl:404:9  */
  assign n12550_o = {n12300_o, n12273_o, n12303_o, n12269_o, n12297_o, n12265_o, n12291_o, n12261_o, n12285_o, n12257_o, n12279_o, n10748_o};
  assign n12553_o = {n9617_o, n9616_o, n9615_o, n9651_o, n12000_o};
  assign n12554_o = {n9621_o, n9518_o, n9655_o, n9511_o, n9510_o, n9654_o, n12001_o};
  assign n12555_o = {n9307_o, 1'b0, 64'b0000000000000000000000000000000000000000000000000000000000000000, n9308_o, 1'b1, n10745_o, n10744_o, n10740_o, n10741_o, n10742_o, n10743_o, c_in, n9311_o, n12004_o};
  assign n12556_o = {n12537_o, n12538_o};
  assign n12557_o = {n12382_o, n12377_o, n12379_o};
  assign n12558_o = {n12440_o, n12434_o, n12428_o, n12422_o, n12416_o, n12410_o, n12404_o, n12398_o, n12390_o, n12392_o};
  reg n12560[61:0] ; // memory
  initial begin
    n12560[61] = 1'b0;
    n12560[60] = 1'b0;
    n12560[59] = 1'b0;
    n12560[58] = 1'b0;
    n12560[57] = 1'b1;
    n12560[56] = 1'b0;
    n12560[55] = 1'b0;
    n12560[54] = 1'b0;
    n12560[53] = 1'b0;
    n12560[52] = 1'b0;
    n12560[51] = 1'b0;
    n12560[50] = 1'b0;
    n12560[49] = 1'b0;
    n12560[48] = 1'b0;
    n12560[47] = 1'b0;
    n12560[46] = 1'b0;
    n12560[45] = 1'b0;
    n12560[44] = 1'b0;
    n12560[43] = 1'b0;
    n12560[42] = 1'b0;
    n12560[41] = 1'b0;
    n12560[40] = 1'b0;
    n12560[39] = 1'b0;
    n12560[38] = 1'b0;
    n12560[37] = 1'b0;
    n12560[36] = 1'b0;
    n12560[35] = 1'b0;
    n12560[34] = 1'b0;
    n12560[33] = 1'b0;
    n12560[32] = 1'b0;
    n12560[31] = 1'b0;
    n12560[30] = 1'b0;
    n12560[29] = 1'b0;
    n12560[28] = 1'b0;
    n12560[27] = 1'b0;
    n12560[26] = 1'b1;
    n12560[25] = 1'b0;
    n12560[24] = 1'b0;
    n12560[23] = 1'b0;
    n12560[22] = 1'b1;
    n12560[21] = 1'b0;
    n12560[20] = 1'b0;
    n12560[19] = 1'b0;
    n12560[18] = 1'b0;
    n12560[17] = 1'b0;
    n12560[16] = 1'b0;
    n12560[15] = 1'b0;
    n12560[14] = 1'b1;
    n12560[13] = 1'b0;
    n12560[12] = 1'b0;
    n12560[11] = 1'b0;
    n12560[10] = 1'b0;
    n12560[9] = 1'b0;
    n12560[8] = 1'b0;
    n12560[7] = 1'b0;
    n12560[6] = 1'b0;
    n12560[5] = 1'b1;
    n12560[4] = 1'b0;
    n12560[3] = 1'b0;
    n12560[2] = 1'b0;
    n12560[1] = 1'b0;
    n12560[0] = 1'b0;
    end
  assign n12561_data = n12560[n10924_o];
  /* execute1.vhdl:166:25  */
  /* execute1.vhdl:166:24  */
  assign n12562_o = cr_in[0];
  /* execute1.vhdl:327:22  */
  assign n12563_o = cr_in[1];
  /* execute1.vhdl:319:20  */
  assign n12564_o = cr_in[2];
  /* execute1.vhdl:318:20  */
  assign n12565_o = cr_in[3];
  /* execute1.vhdl:317:21  */
  assign n12566_o = cr_in[4];
  /* execute1.vhdl:311:22  */
  assign n12567_o = cr_in[5];
  /* execute1.vhdl:303:22  */
  assign n12568_o = cr_in[6];
  /* execute1.vhdl:296:23  */
  assign n12569_o = cr_in[7];
  /* execute1.vhdl:284:23  */
  assign n12570_o = cr_in[8];
  /* execute1.vhdl:274:26  */
  assign n12571_o = cr_in[9];
  /* execute1.vhdl:273:23  */
  assign n12572_o = cr_in[10];
  /* execute1.vhdl:56:9  */
  assign n12573_o = cr_in[11];
  /* execute1.vhdl:55:9  */
  assign n12574_o = cr_in[12];
  /* execute1.vhdl:47:9  */
  assign n12575_o = cr_in[13];
  /* execute1.vhdl:46:9  */
  assign n12576_o = cr_in[14];
  /* execute1.vhdl:44:9  */
  assign n12577_o = cr_in[15];
  /* execute1.vhdl:42:9  */
  assign n12578_o = cr_in[16];
  /* execute1.vhdl:41:9  */
  assign n12579_o = cr_in[17];
  /* execute1.vhdl:40:9  */
  assign n12580_o = cr_in[18];
  /* execute1.vhdl:38:9  */
  assign n12581_o = cr_in[19];
  /* execute1.vhdl:37:9  */
  assign n12582_o = cr_in[20];
  /* execute1.vhdl:27:9  */
  assign n12583_o = cr_in[21];
  assign n12584_o = cr_in[22];
  assign n12585_o = cr_in[23];
  assign n12586_o = cr_in[24];
  assign n12587_o = cr_in[25];
  assign n12588_o = cr_in[26];
  assign n12589_o = cr_in[27];
  assign n12590_o = cr_in[28];
  assign n12591_o = cr_in[29];
  assign n12592_o = cr_in[30];
  assign n12593_o = cr_in[31];
  /* execute1.vhdl:581:25  */
  assign n12594_o = n9843_o[1:0];
  /* execute1.vhdl:581:25  */
  always @*
    case (n12594_o)
      2'b00: n12595_o = n12562_o;
      2'b01: n12595_o = n12563_o;
      2'b10: n12595_o = n12564_o;
      2'b11: n12595_o = n12565_o;
    endcase
  /* execute1.vhdl:581:25  */
  assign n12596_o = n9843_o[1:0];
  /* execute1.vhdl:581:25  */
  always @*
    case (n12596_o)
      2'b00: n12597_o = n12566_o;
      2'b01: n12597_o = n12567_o;
      2'b10: n12597_o = n12568_o;
      2'b11: n12597_o = n12569_o;
    endcase
  /* execute1.vhdl:581:25  */
  assign n12598_o = n9843_o[1:0];
  /* execute1.vhdl:581:25  */
  always @*
    case (n12598_o)
      2'b00: n12599_o = n12570_o;
      2'b01: n12599_o = n12571_o;
      2'b10: n12599_o = n12572_o;
      2'b11: n12599_o = n12573_o;
    endcase
  /* execute1.vhdl:581:25  */
  assign n12600_o = n9843_o[1:0];
  /* execute1.vhdl:581:25  */
  always @*
    case (n12600_o)
      2'b00: n12601_o = n12574_o;
      2'b01: n12601_o = n12575_o;
      2'b10: n12601_o = n12576_o;
      2'b11: n12601_o = n12577_o;
    endcase
  /* execute1.vhdl:581:25  */
  assign n12602_o = n9843_o[1:0];
  /* execute1.vhdl:581:25  */
  always @*
    case (n12602_o)
      2'b00: n12603_o = n12578_o;
      2'b01: n12603_o = n12579_o;
      2'b10: n12603_o = n12580_o;
      2'b11: n12603_o = n12581_o;
    endcase
  /* execute1.vhdl:581:25  */
  assign n12604_o = n9843_o[1:0];
  /* execute1.vhdl:581:25  */
  always @*
    case (n12604_o)
      2'b00: n12605_o = n12582_o;
      2'b01: n12605_o = n12583_o;
      2'b10: n12605_o = n12584_o;
      2'b11: n12605_o = n12585_o;
    endcase
  /* execute1.vhdl:581:25  */
  assign n12606_o = n9843_o[1:0];
  /* execute1.vhdl:581:25  */
  always @*
    case (n12606_o)
      2'b00: n12607_o = n12586_o;
      2'b01: n12607_o = n12587_o;
      2'b10: n12607_o = n12588_o;
      2'b11: n12607_o = n12589_o;
    endcase
  /* execute1.vhdl:581:25  */
  assign n12608_o = n9843_o[1:0];
  /* execute1.vhdl:581:25  */
  always @*
    case (n12608_o)
      2'b00: n12609_o = n12590_o;
      2'b01: n12609_o = n12591_o;
      2'b10: n12609_o = n12592_o;
      2'b11: n12609_o = n12593_o;
    endcase
  /* execute1.vhdl:581:25  */
  assign n12610_o = n9843_o[3:2];
  /* execute1.vhdl:581:25  */
  always @*
    case (n12610_o)
      2'b00: n12611_o = n12595_o;
      2'b01: n12611_o = n12597_o;
      2'b10: n12611_o = n12599_o;
      2'b11: n12611_o = n12601_o;
    endcase
  /* execute1.vhdl:581:25  */
  assign n12612_o = n9843_o[3:2];
  /* execute1.vhdl:581:25  */
  always @*
    case (n12612_o)
      2'b00: n12613_o = n12603_o;
      2'b01: n12613_o = n12605_o;
      2'b10: n12613_o = n12607_o;
      2'b11: n12613_o = n12609_o;
    endcase
  /* execute1.vhdl:581:25  */
  assign n12614_o = n9843_o[4];
  /* execute1.vhdl:581:25  */
  assign n12615_o = n12614_o ? n12613_o : n12611_o;
  /* execute1.vhdl:581:25  */
  assign n12616_o = cr_in[0];
  /* execute1.vhdl:581:28  */
  assign n12617_o = cr_in[1];
  assign n12618_o = cr_in[2];
  assign n12619_o = cr_in[3];
  assign n12620_o = cr_in[4];
  assign n12621_o = cr_in[5];
  assign n12622_o = cr_in[6];
  assign n12623_o = cr_in[7];
  assign n12624_o = cr_in[8];
  assign n12625_o = cr_in[9];
  assign n12626_o = cr_in[10];
  assign n12627_o = cr_in[11];
  assign n12628_o = cr_in[12];
  assign n12629_o = cr_in[13];
  assign n12630_o = cr_in[14];
  assign n12631_o = cr_in[15];
  assign n12632_o = cr_in[16];
  assign n12633_o = cr_in[17];
  assign n12634_o = cr_in[18];
  assign n12635_o = cr_in[19];
  /* execute1.vhdl:913:9  */
  assign n12636_o = cr_in[20];
  assign n12637_o = cr_in[21];
  assign n12638_o = cr_in[22];
  /* execute1.vhdl:913:9  */
  assign n12639_o = cr_in[23];
  assign n12640_o = cr_in[24];
  assign n12641_o = cr_in[25];
  /* execute1.vhdl:913:9  */
  assign n12642_o = cr_in[26];
  assign n12643_o = cr_in[27];
  assign n12644_o = cr_in[28];
  /* execute1.vhdl:913:9  */
  assign n12645_o = cr_in[29];
  assign n12646_o = cr_in[30];
  assign n12647_o = cr_in[31];
  /* execute1.vhdl:626:25  */
  assign n12648_o = n10072_o[1:0];
  /* execute1.vhdl:626:25  */
  always @*
    case (n12648_o)
      2'b00: n12649_o = n12616_o;
      2'b01: n12649_o = n12617_o;
      2'b10: n12649_o = n12618_o;
      2'b11: n12649_o = n12619_o;
    endcase
  /* execute1.vhdl:626:25  */
  assign n12650_o = n10072_o[1:0];
  /* execute1.vhdl:626:25  */
  always @*
    case (n12650_o)
      2'b00: n12651_o = n12620_o;
      2'b01: n12651_o = n12621_o;
      2'b10: n12651_o = n12622_o;
      2'b11: n12651_o = n12623_o;
    endcase
  /* execute1.vhdl:626:25  */
  assign n12652_o = n10072_o[1:0];
  /* execute1.vhdl:626:25  */
  always @*
    case (n12652_o)
      2'b00: n12653_o = n12624_o;
      2'b01: n12653_o = n12625_o;
      2'b10: n12653_o = n12626_o;
      2'b11: n12653_o = n12627_o;
    endcase
  /* execute1.vhdl:626:25  */
  assign n12654_o = n10072_o[1:0];
  /* execute1.vhdl:626:25  */
  always @*
    case (n12654_o)
      2'b00: n12655_o = n12628_o;
      2'b01: n12655_o = n12629_o;
      2'b10: n12655_o = n12630_o;
      2'b11: n12655_o = n12631_o;
    endcase
  /* execute1.vhdl:626:25  */
  assign n12656_o = n10072_o[1:0];
  /* execute1.vhdl:626:25  */
  always @*
    case (n12656_o)
      2'b00: n12657_o = n12632_o;
      2'b01: n12657_o = n12633_o;
      2'b10: n12657_o = n12634_o;
      2'b11: n12657_o = n12635_o;
    endcase
  /* execute1.vhdl:626:25  */
  assign n12658_o = n10072_o[1:0];
  /* execute1.vhdl:626:25  */
  always @*
    case (n12658_o)
      2'b00: n12659_o = n12636_o;
      2'b01: n12659_o = n12637_o;
      2'b10: n12659_o = n12638_o;
      2'b11: n12659_o = n12639_o;
    endcase
  /* execute1.vhdl:626:25  */
  assign n12660_o = n10072_o[1:0];
  /* execute1.vhdl:626:25  */
  always @*
    case (n12660_o)
      2'b00: n12661_o = n12640_o;
      2'b01: n12661_o = n12641_o;
      2'b10: n12661_o = n12642_o;
      2'b11: n12661_o = n12643_o;
    endcase
  /* execute1.vhdl:626:25  */
  assign n12662_o = n10072_o[1:0];
  /* execute1.vhdl:626:25  */
  always @*
    case (n12662_o)
      2'b00: n12663_o = n12644_o;
      2'b01: n12663_o = n12645_o;
      2'b10: n12663_o = n12646_o;
      2'b11: n12663_o = n12647_o;
    endcase
  /* execute1.vhdl:626:25  */
  assign n12664_o = n10072_o[3:2];
  /* execute1.vhdl:626:25  */
  always @*
    case (n12664_o)
      2'b00: n12665_o = n12649_o;
      2'b01: n12665_o = n12651_o;
      2'b10: n12665_o = n12653_o;
      2'b11: n12665_o = n12655_o;
    endcase
  /* execute1.vhdl:626:25  */
  assign n12666_o = n10072_o[3:2];
  /* execute1.vhdl:626:25  */
  always @*
    case (n12666_o)
      2'b00: n12667_o = n12657_o;
      2'b01: n12667_o = n12659_o;
      2'b10: n12667_o = n12661_o;
      2'b11: n12667_o = n12663_o;
    endcase
  /* execute1.vhdl:626:25  */
  assign n12668_o = n10072_o[4];
  /* execute1.vhdl:626:25  */
  assign n12669_o = n12668_o ? n12667_o : n12665_o;
  /* execute1.vhdl:626:25  */
  assign n12670_o = cr_in[0];
  /* execute1.vhdl:626:29  */
  assign n12671_o = cr_in[1];
  assign n12672_o = cr_in[2];
  assign n12673_o = cr_in[3];
  assign n12674_o = cr_in[4];
  /* execute1.vhdl:913:9  */
  assign n12675_o = cr_in[5];
  assign n12676_o = cr_in[6];
  assign n12677_o = cr_in[7];
  /* execute1.vhdl:913:9  */
  assign n12678_o = cr_in[8];
  assign n12679_o = cr_in[9];
  assign n12680_o = cr_in[10];
  /* execute1.vhdl:913:9  */
  assign n12681_o = cr_in[11];
  assign n12682_o = cr_in[12];
  assign n12683_o = cr_in[13];
  /* execute1.vhdl:913:9  */
  assign n12684_o = cr_in[14];
  assign n12685_o = cr_in[15];
  assign n12686_o = cr_in[16];
  /* execute1.vhdl:913:9  */
  assign n12687_o = cr_in[17];
  assign n12688_o = cr_in[18];
  assign n12689_o = cr_in[19];
  assign n12690_o = cr_in[20];
  /* execute1.vhdl:913:9  */
  assign n12691_o = cr_in[21];
  /* execute1.vhdl:913:9  */
  assign n12692_o = cr_in[22];
  /* execute1.vhdl:913:9  */
  assign n12693_o = cr_in[23];
  /* execute1.vhdl:913:9  */
  assign n12694_o = cr_in[24];
  /* execute1.vhdl:913:9  */
  assign n12695_o = cr_in[25];
  /* execute1.vhdl:913:9  */
  assign n12696_o = cr_in[26];
  assign n12697_o = cr_in[27];
  /* execute1.vhdl:913:9  */
  assign n12698_o = cr_in[28];
  assign n12699_o = cr_in[29];
  assign n12700_o = cr_in[30];
  /* execute1.vhdl:916:13  */
  assign n12701_o = cr_in[31];
  /* execute1.vhdl:628:28  */
  assign n12702_o = n10078_o[1:0];
  /* execute1.vhdl:628:28  */
  always @*
    case (n12702_o)
      2'b00: n12703_o = n12670_o;
      2'b01: n12703_o = n12671_o;
      2'b10: n12703_o = n12672_o;
      2'b11: n12703_o = n12673_o;
    endcase
  /* execute1.vhdl:628:28  */
  assign n12704_o = n10078_o[1:0];
  /* execute1.vhdl:628:28  */
  always @*
    case (n12704_o)
      2'b00: n12705_o = n12674_o;
      2'b01: n12705_o = n12675_o;
      2'b10: n12705_o = n12676_o;
      2'b11: n12705_o = n12677_o;
    endcase
  /* execute1.vhdl:628:28  */
  assign n12706_o = n10078_o[1:0];
  /* execute1.vhdl:628:28  */
  always @*
    case (n12706_o)
      2'b00: n12707_o = n12678_o;
      2'b01: n12707_o = n12679_o;
      2'b10: n12707_o = n12680_o;
      2'b11: n12707_o = n12681_o;
    endcase
  /* execute1.vhdl:628:28  */
  assign n12708_o = n10078_o[1:0];
  /* execute1.vhdl:628:28  */
  always @*
    case (n12708_o)
      2'b00: n12709_o = n12682_o;
      2'b01: n12709_o = n12683_o;
      2'b10: n12709_o = n12684_o;
      2'b11: n12709_o = n12685_o;
    endcase
  /* execute1.vhdl:628:28  */
  assign n12710_o = n10078_o[1:0];
  /* execute1.vhdl:628:28  */
  always @*
    case (n12710_o)
      2'b00: n12711_o = n12686_o;
      2'b01: n12711_o = n12687_o;
      2'b10: n12711_o = n12688_o;
      2'b11: n12711_o = n12689_o;
    endcase
  /* execute1.vhdl:628:28  */
  assign n12712_o = n10078_o[1:0];
  /* execute1.vhdl:628:28  */
  always @*
    case (n12712_o)
      2'b00: n12713_o = n12690_o;
      2'b01: n12713_o = n12691_o;
      2'b10: n12713_o = n12692_o;
      2'b11: n12713_o = n12693_o;
    endcase
  /* execute1.vhdl:628:28  */
  assign n12714_o = n10078_o[1:0];
  /* execute1.vhdl:628:28  */
  always @*
    case (n12714_o)
      2'b00: n12715_o = n12694_o;
      2'b01: n12715_o = n12695_o;
      2'b10: n12715_o = n12696_o;
      2'b11: n12715_o = n12697_o;
    endcase
  /* execute1.vhdl:628:28  */
  assign n12716_o = n10078_o[1:0];
  /* execute1.vhdl:628:28  */
  always @*
    case (n12716_o)
      2'b00: n12717_o = n12698_o;
      2'b01: n12717_o = n12699_o;
      2'b10: n12717_o = n12700_o;
      2'b11: n12717_o = n12701_o;
    endcase
  /* execute1.vhdl:628:28  */
  assign n12718_o = n10078_o[3:2];
  /* execute1.vhdl:628:28  */
  always @*
    case (n12718_o)
      2'b00: n12719_o = n12703_o;
      2'b01: n12719_o = n12705_o;
      2'b10: n12719_o = n12707_o;
      2'b11: n12719_o = n12709_o;
    endcase
  /* execute1.vhdl:628:28  */
  assign n12720_o = n10078_o[3:2];
  /* execute1.vhdl:628:28  */
  always @*
    case (n12720_o)
      2'b00: n12721_o = n12711_o;
      2'b01: n12721_o = n12713_o;
      2'b10: n12721_o = n12715_o;
      2'b11: n12721_o = n12717_o;
    endcase
  /* execute1.vhdl:628:28  */
  assign n12722_o = n10078_o[4];
  /* execute1.vhdl:628:28  */
  assign n12723_o = n12722_o ? n12721_o : n12719_o;
  /* execute1.vhdl:628:28  */
  assign n12724_o = cr_in[3:0];
  /* execute1.vhdl:628:32  */
  assign n12725_o = cr_in[7:4];
  assign n12726_o = cr_in[11:8];
  /* common.vhdl:112:14  */
  assign n12727_o = cr_in[15:12];
  /* common.vhdl:112:14  */
  assign n12728_o = cr_in[19:16];
  assign n12729_o = cr_in[23:20];
  /* common.vhdl:112:14  */
  assign n12730_o = cr_in[27:24];
  /* common.vhdl:708:16  */
  assign n12731_o = cr_in[31:28];
  /* execute1.vhdl:699:36  */
  assign n12732_o = n10342_o[1:0];
  /* execute1.vhdl:699:36  */
  always @*
    case (n12732_o)
      2'b00: n12733_o = n12724_o;
      2'b01: n12733_o = n12725_o;
      2'b10: n12733_o = n12726_o;
      2'b11: n12733_o = n12727_o;
    endcase
  /* execute1.vhdl:699:36  */
  assign n12734_o = n10342_o[1:0];
  /* execute1.vhdl:699:36  */
  always @*
    case (n12734_o)
      2'b00: n12735_o = n12728_o;
      2'b01: n12735_o = n12729_o;
      2'b10: n12735_o = n12730_o;
      2'b11: n12735_o = n12731_o;
    endcase
  /* execute1.vhdl:699:36  */
  assign n12736_o = n10342_o[2];
  /* execute1.vhdl:699:36  */
  assign n12737_o = n12736_o ? n12735_o : n12733_o;
  /* execute1.vhdl:699:36  */
  assign n12738_o = cr_in[0];
  /* execute1.vhdl:699:36  */
  assign n12739_o = cr_in[1];
  /* common.vhdl:31:14  */
  assign n12740_o = cr_in[2];
  assign n12741_o = cr_in[3];
  /* common.vhdl:31:14  */
  assign n12742_o = cr_in[4];
  /* common.vhdl:112:14  */
  assign n12743_o = cr_in[5];
  /* common.vhdl:112:14  */
  assign n12744_o = cr_in[6];
  assign n12745_o = cr_in[7];
  /* common.vhdl:112:14  */
  assign n12746_o = cr_in[8];
  assign n12747_o = cr_in[9];
  /* execute1.vhdl:1017:51  */
  assign n12748_o = cr_in[10];
  assign n12749_o = cr_in[11];
  assign n12750_o = cr_in[12];
  assign n12751_o = cr_in[13];
  assign n12752_o = cr_in[14];
  assign n12753_o = cr_in[15];
  /* ppc_fx_insns.vhdl:823:26  */
  assign n12754_o = cr_in[16];
  assign n12755_o = cr_in[17];
  /* ppc_fx_insns.vhdl:822:26  */
  assign n12756_o = cr_in[18];
  assign n12757_o = cr_in[19];
  /* ppc_fx_insns.vhdl:821:26  */
  assign n12758_o = cr_in[20];
  assign n12759_o = cr_in[21];
  /* ppc_fx_insns.vhdl:820:26  */
  assign n12760_o = cr_in[22];
  assign n12761_o = cr_in[23];
  /* ppc_fx_insns.vhdl:819:26  */
  assign n12762_o = cr_in[24];
  assign n12763_o = cr_in[25];
  /* ppc_fx_insns.vhdl:98:18  */
  assign n12764_o = cr_in[26];
  /* ppc_fx_insns.vhdl:98:18  */
  assign n12765_o = cr_in[27];
  assign n12766_o = cr_in[28];
  /* ppc_fx_insns.vhdl:98:18  */
  assign n12767_o = cr_in[29];
  /* insn_helpers.vhdl:30:14  */
  assign n12768_o = cr_in[30];
  /* insn_helpers.vhdl:30:14  */
  assign n12769_o = cr_in[31];
  /* execute1.vhdl:708:41  */
  assign n12770_o = n10376_o[1:0];
  /* execute1.vhdl:708:41  */
  always @*
    case (n12770_o)
      2'b00: n12771_o = n12738_o;
      2'b01: n12771_o = n12739_o;
      2'b10: n12771_o = n12740_o;
      2'b11: n12771_o = n12741_o;
    endcase
  /* execute1.vhdl:708:41  */
  assign n12772_o = n10376_o[1:0];
  /* execute1.vhdl:708:41  */
  always @*
    case (n12772_o)
      2'b00: n12773_o = n12742_o;
      2'b01: n12773_o = n12743_o;
      2'b10: n12773_o = n12744_o;
      2'b11: n12773_o = n12745_o;
    endcase
  /* execute1.vhdl:708:41  */
  assign n12774_o = n10376_o[1:0];
  /* execute1.vhdl:708:41  */
  always @*
    case (n12774_o)
      2'b00: n12775_o = n12746_o;
      2'b01: n12775_o = n12747_o;
      2'b10: n12775_o = n12748_o;
      2'b11: n12775_o = n12749_o;
    endcase
  /* execute1.vhdl:708:41  */
  assign n12776_o = n10376_o[1:0];
  /* execute1.vhdl:708:41  */
  always @*
    case (n12776_o)
      2'b00: n12777_o = n12750_o;
      2'b01: n12777_o = n12751_o;
      2'b10: n12777_o = n12752_o;
      2'b11: n12777_o = n12753_o;
    endcase
  /* execute1.vhdl:708:41  */
  assign n12778_o = n10376_o[1:0];
  /* execute1.vhdl:708:41  */
  always @*
    case (n12778_o)
      2'b00: n12779_o = n12754_o;
      2'b01: n12779_o = n12755_o;
      2'b10: n12779_o = n12756_o;
      2'b11: n12779_o = n12757_o;
    endcase
  /* execute1.vhdl:708:41  */
  assign n12780_o = n10376_o[1:0];
  /* execute1.vhdl:708:41  */
  always @*
    case (n12780_o)
      2'b00: n12781_o = n12758_o;
      2'b01: n12781_o = n12759_o;
      2'b10: n12781_o = n12760_o;
      2'b11: n12781_o = n12761_o;
    endcase
  /* execute1.vhdl:708:41  */
  assign n12782_o = n10376_o[1:0];
  /* execute1.vhdl:708:41  */
  always @*
    case (n12782_o)
      2'b00: n12783_o = n12762_o;
      2'b01: n12783_o = n12763_o;
      2'b10: n12783_o = n12764_o;
      2'b11: n12783_o = n12765_o;
    endcase
  /* execute1.vhdl:708:41  */
  assign n12784_o = n10376_o[1:0];
  /* execute1.vhdl:708:41  */
  always @*
    case (n12784_o)
      2'b00: n12785_o = n12766_o;
      2'b01: n12785_o = n12767_o;
      2'b10: n12785_o = n12768_o;
      2'b11: n12785_o = n12769_o;
    endcase
  /* execute1.vhdl:708:41  */
  assign n12786_o = n10376_o[3:2];
  /* execute1.vhdl:708:41  */
  always @*
    case (n12786_o)
      2'b00: n12787_o = n12771_o;
      2'b01: n12787_o = n12773_o;
      2'b10: n12787_o = n12775_o;
      2'b11: n12787_o = n12777_o;
    endcase
  /* execute1.vhdl:708:41  */
  assign n12788_o = n10376_o[3:2];
  /* execute1.vhdl:708:41  */
  always @*
    case (n12788_o)
      2'b00: n12789_o = n12779_o;
      2'b01: n12789_o = n12781_o;
      2'b10: n12789_o = n12783_o;
      2'b11: n12789_o = n12785_o;
    endcase
  /* execute1.vhdl:708:41  */
  assign n12790_o = n10376_o[4];
  /* execute1.vhdl:708:41  */
  assign n12791_o = n12790_o ? n12789_o : n12787_o;
  /* execute1.vhdl:708:41  */
  assign n12792_o = cr_in[0];
  /* execute1.vhdl:708:42  */
  assign n12793_o = cr_in[1];
  assign n12794_o = cr_in[2];
  /* execute1.vhdl:822:9  */
  assign n12795_o = cr_in[3];
  assign n12796_o = cr_in[4];
  assign n12797_o = cr_in[5];
  /* execute1.vhdl:822:9  */
  assign n12798_o = cr_in[6];
  assign n12799_o = cr_in[7];
  assign n12800_o = cr_in[8];
  /* execute1.vhdl:163:14  */
  assign n12801_o = cr_in[9];
  /* execute1.vhdl:163:14  */
  assign n12802_o = cr_in[10];
  assign n12803_o = cr_in[11];
  /* execute1.vhdl:163:14  */
  assign n12804_o = cr_in[12];
  assign n12805_o = cr_in[13];
  assign n12806_o = cr_in[14];
  assign n12807_o = cr_in[15];
  /* execute1.vhdl:822:9  */
  assign n12808_o = cr_in[16];
  assign n12809_o = cr_in[17];
  /* execute1.vhdl:823:29  */
  assign n12810_o = cr_in[18];
  /* execute1.vhdl:823:27  */
  assign n12811_o = cr_in[19];
  assign n12812_o = cr_in[20];
  assign n12813_o = cr_in[21];
  assign n12814_o = cr_in[22];
  assign n12815_o = cr_in[23];
  assign n12816_o = cr_in[24];
  assign n12817_o = cr_in[25];
  assign n12818_o = cr_in[26];
  assign n12819_o = cr_in[27];
  assign n12820_o = cr_in[28];
  assign n12821_o = cr_in[29];
  assign n12822_o = cr_in[30];
  assign n12823_o = cr_in[31];
  /* execute1.vhdl:708:56  */
  assign n12824_o = n10381_o[1:0];
  /* execute1.vhdl:708:56  */
  always @*
    case (n12824_o)
      2'b00: n12825_o = n12792_o;
      2'b01: n12825_o = n12793_o;
      2'b10: n12825_o = n12794_o;
      2'b11: n12825_o = n12795_o;
    endcase
  /* execute1.vhdl:708:56  */
  assign n12826_o = n10381_o[1:0];
  /* execute1.vhdl:708:56  */
  always @*
    case (n12826_o)
      2'b00: n12827_o = n12796_o;
      2'b01: n12827_o = n12797_o;
      2'b10: n12827_o = n12798_o;
      2'b11: n12827_o = n12799_o;
    endcase
  /* execute1.vhdl:708:56  */
  assign n12828_o = n10381_o[1:0];
  /* execute1.vhdl:708:56  */
  always @*
    case (n12828_o)
      2'b00: n12829_o = n12800_o;
      2'b01: n12829_o = n12801_o;
      2'b10: n12829_o = n12802_o;
      2'b11: n12829_o = n12803_o;
    endcase
  /* execute1.vhdl:708:56  */
  assign n12830_o = n10381_o[1:0];
  /* execute1.vhdl:708:56  */
  always @*
    case (n12830_o)
      2'b00: n12831_o = n12804_o;
      2'b01: n12831_o = n12805_o;
      2'b10: n12831_o = n12806_o;
      2'b11: n12831_o = n12807_o;
    endcase
  /* execute1.vhdl:708:56  */
  assign n12832_o = n10381_o[1:0];
  /* execute1.vhdl:708:56  */
  always @*
    case (n12832_o)
      2'b00: n12833_o = n12808_o;
      2'b01: n12833_o = n12809_o;
      2'b10: n12833_o = n12810_o;
      2'b11: n12833_o = n12811_o;
    endcase
  /* execute1.vhdl:708:56  */
  assign n12834_o = n10381_o[1:0];
  /* execute1.vhdl:708:56  */
  always @*
    case (n12834_o)
      2'b00: n12835_o = n12812_o;
      2'b01: n12835_o = n12813_o;
      2'b10: n12835_o = n12814_o;
      2'b11: n12835_o = n12815_o;
    endcase
  /* execute1.vhdl:708:56  */
  assign n12836_o = n10381_o[1:0];
  /* execute1.vhdl:708:56  */
  always @*
    case (n12836_o)
      2'b00: n12837_o = n12816_o;
      2'b01: n12837_o = n12817_o;
      2'b10: n12837_o = n12818_o;
      2'b11: n12837_o = n12819_o;
    endcase
  /* execute1.vhdl:708:56  */
  assign n12838_o = n10381_o[1:0];
  /* execute1.vhdl:708:56  */
  always @*
    case (n12838_o)
      2'b00: n12839_o = n12820_o;
      2'b01: n12839_o = n12821_o;
      2'b10: n12839_o = n12822_o;
      2'b11: n12839_o = n12823_o;
    endcase
  /* execute1.vhdl:708:56  */
  assign n12840_o = n10381_o[3:2];
  /* execute1.vhdl:708:56  */
  always @*
    case (n12840_o)
      2'b00: n12841_o = n12825_o;
      2'b01: n12841_o = n12827_o;
      2'b10: n12841_o = n12829_o;
      2'b11: n12841_o = n12831_o;
    endcase
  /* execute1.vhdl:708:56  */
  assign n12842_o = n10381_o[3:2];
  /* execute1.vhdl:708:56  */
  always @*
    case (n12842_o)
      2'b00: n12843_o = n12833_o;
      2'b01: n12843_o = n12835_o;
      2'b10: n12843_o = n12837_o;
      2'b11: n12843_o = n12839_o;
    endcase
  /* execute1.vhdl:708:56  */
  assign n12844_o = n10381_o[4];
  /* execute1.vhdl:708:56  */
  assign n12845_o = n12844_o ? n12843_o : n12841_o;
  /* execute1.vhdl:708:56  */
  assign n12846_o = n9139_o[343];
  /* execute1.vhdl:708:57  */
  assign n12847_o = n9139_o[344];
  assign n12848_o = n9139_o[345];
  /* execute1.vhdl:751:18  */
  assign n12849_o = n9139_o[346];
  assign n12850_o = n9139_o[347];
  /* execute1.vhdl:750:18  */
  assign n12851_o = n9139_o[348];
  assign n12852_o = n9139_o[349];
  /* execute1.vhdl:749:18  */
  assign n12853_o = n9139_o[350];
  assign n12854_o = n9139_o[351];
  /* execute1.vhdl:748:18  */
  assign n12855_o = n9139_o[352];
  assign n12856_o = n9139_o[353];
  /* execute1.vhdl:747:22  */
  assign n12857_o = n9139_o[354];
  assign n12858_o = n9139_o[355];
  /* execute1.vhdl:747:18  */
  assign n12859_o = n9139_o[356];
  assign n12860_o = n9139_o[357];
  /* execute1.vhdl:746:18  */
  assign n12861_o = n9139_o[358];
  assign n12862_o = n9139_o[359];
  assign n12863_o = n9139_o[360];
  assign n12864_o = n9139_o[361];
  assign n12865_o = n9139_o[362];
  /* execute1.vhdl:727:9  */
  assign n12866_o = n9139_o[363];
  /* crhelpers.vhdl:12:14  */
  assign n12867_o = n9139_o[364];
  /* crhelpers.vhdl:12:14  */
  assign n12868_o = n9139_o[365];
  assign n12869_o = n9139_o[366];
  /* crhelpers.vhdl:12:14  */
  assign n12870_o = n9139_o[367];
  /* execute1.vhdl:728:13  */
  assign n12871_o = n9139_o[368];
  /* crhelpers.vhdl:12:14  */
  assign n12872_o = n9139_o[369];
  /* crhelpers.vhdl:12:14  */
  assign n12873_o = n9139_o[370];
  assign n12874_o = n9139_o[371];
  /* crhelpers.vhdl:12:14  */
  assign n12875_o = n9139_o[372];
  /* crhelpers.vhdl:30:9  */
  assign n12876_o = n9139_o[373];
  assign n12877_o = n9139_o[374];
  /* execute1.vhdl:709:42  */
  assign n12878_o = n10391_o[1:0];
  /* execute1.vhdl:709:42  */
  always @*
    case (n12878_o)
      2'b00: n12879_o = n12846_o;
      2'b01: n12879_o = n12847_o;
      2'b10: n12879_o = n12848_o;
      2'b11: n12879_o = n12849_o;
    endcase
  /* execute1.vhdl:709:42  */
  assign n12880_o = n10391_o[1:0];
  /* execute1.vhdl:709:42  */
  always @*
    case (n12880_o)
      2'b00: n12881_o = n12850_o;
      2'b01: n12881_o = n12851_o;
      2'b10: n12881_o = n12852_o;
      2'b11: n12881_o = n12853_o;
    endcase
  /* execute1.vhdl:709:42  */
  assign n12882_o = n10391_o[1:0];
  /* execute1.vhdl:709:42  */
  always @*
    case (n12882_o)
      2'b00: n12883_o = n12854_o;
      2'b01: n12883_o = n12855_o;
      2'b10: n12883_o = n12856_o;
      2'b11: n12883_o = n12857_o;
    endcase
  /* execute1.vhdl:709:42  */
  assign n12884_o = n10391_o[1:0];
  /* execute1.vhdl:709:42  */
  always @*
    case (n12884_o)
      2'b00: n12885_o = n12858_o;
      2'b01: n12885_o = n12859_o;
      2'b10: n12885_o = n12860_o;
      2'b11: n12885_o = n12861_o;
    endcase
  /* execute1.vhdl:709:42  */
  assign n12886_o = n10391_o[1:0];
  /* execute1.vhdl:709:42  */
  always @*
    case (n12886_o)
      2'b00: n12887_o = n12862_o;
      2'b01: n12887_o = n12863_o;
      2'b10: n12887_o = n12864_o;
      2'b11: n12887_o = n12865_o;
    endcase
  /* execute1.vhdl:709:42  */
  assign n12888_o = n10391_o[1:0];
  /* execute1.vhdl:709:42  */
  always @*
    case (n12888_o)
      2'b00: n12889_o = n12866_o;
      2'b01: n12889_o = n12867_o;
      2'b10: n12889_o = n12868_o;
      2'b11: n12889_o = n12869_o;
    endcase
  /* execute1.vhdl:709:42  */
  assign n12890_o = n10391_o[1:0];
  /* execute1.vhdl:709:42  */
  always @*
    case (n12890_o)
      2'b00: n12891_o = n12870_o;
      2'b01: n12891_o = n12871_o;
      2'b10: n12891_o = n12872_o;
      2'b11: n12891_o = n12873_o;
    endcase
  /* execute1.vhdl:709:42  */
  assign n12892_o = n10391_o[1:0];
  /* execute1.vhdl:709:42  */
  always @*
    case (n12892_o)
      2'b00: n12893_o = n12874_o;
      2'b01: n12893_o = n12875_o;
      2'b10: n12893_o = n12876_o;
      2'b11: n12893_o = n12877_o;
    endcase
  /* execute1.vhdl:709:42  */
  assign n12894_o = n10391_o[3:2];
  /* execute1.vhdl:709:42  */
  always @*
    case (n12894_o)
      2'b00: n12895_o = n12879_o;
      2'b01: n12895_o = n12881_o;
      2'b10: n12895_o = n12883_o;
      2'b11: n12895_o = n12885_o;
    endcase
  /* execute1.vhdl:709:42  */
  assign n12896_o = n10391_o[3:2];
  /* execute1.vhdl:709:42  */
  always @*
    case (n12896_o)
      2'b00: n12897_o = n12887_o;
      2'b01: n12897_o = n12889_o;
      2'b10: n12897_o = n12891_o;
      2'b11: n12897_o = n12893_o;
    endcase
  /* execute1.vhdl:709:42  */
  assign n12898_o = n10391_o[4];
  /* execute1.vhdl:709:42  */
  assign n12899_o = n12898_o ? n12897_o : n12895_o;
  /* execute1.vhdl:709:42  */
  assign n12900_o = cr_in[3:0];
  /* execute1.vhdl:709:45  */
  assign n12901_o = cr_in[7:4];
  /* execute1.vhdl:683:9  */
  assign n12902_o = cr_in[11:8];
  /* execute1.vhdl:683:9  */
  assign n12903_o = cr_in[15:12];
  /* execute1.vhdl:683:9  */
  assign n12904_o = cr_in[19:16];
  /* execute1.vhdl:683:9  */
  assign n12905_o = cr_in[23:20];
  /* execute1.vhdl:683:9  */
  assign n12906_o = cr_in[27:24];
  /* execute1.vhdl:683:9  */
  assign n12907_o = cr_in[31:28];
  /* execute1.vhdl:720:36  */
  assign n12908_o = n10432_o[1:0];
  /* execute1.vhdl:720:36  */
  always @*
    case (n12908_o)
      2'b00: n12909_o = n12900_o;
      2'b01: n12909_o = n12901_o;
      2'b10: n12909_o = n12902_o;
      2'b11: n12909_o = n12903_o;
    endcase
  /* execute1.vhdl:720:36  */
  assign n12910_o = n10432_o[1:0];
  /* execute1.vhdl:720:36  */
  always @*
    case (n12910_o)
      2'b00: n12911_o = n12904_o;
      2'b01: n12911_o = n12905_o;
      2'b10: n12911_o = n12906_o;
      2'b11: n12911_o = n12907_o;
    endcase
  /* execute1.vhdl:720:36  */
  assign n12912_o = n10432_o[2];
  /* execute1.vhdl:720:36  */
  assign n12913_o = n12912_o ? n12911_o : n12909_o;
  /* execute1.vhdl:720:36  */
  assign n12914_o = cr_in[0];
  /* execute1.vhdl:720:36  */
  assign n12915_o = cr_in[1];
  /* execute1.vhdl:696:17  */
  assign n12916_o = cr_in[2];
  /* execute1.vhdl:696:17  */
  assign n12917_o = cr_in[3];
  /* execute1.vhdl:696:17  */
  assign n12918_o = cr_in[4];
  /* execute1.vhdl:696:17  */
  assign n12919_o = cr_in[5];
  /* execute1.vhdl:696:17  */
  assign n12920_o = cr_in[6];
  /* execute1.vhdl:696:17  */
  assign n12921_o = cr_in[7];
  /* execute1.vhdl:696:17  */
  assign n12922_o = cr_in[8];
  /* execute1.vhdl:696:17  */
  assign n12923_o = cr_in[9];
  /* execute1.vhdl:720:39  */
  assign n12924_o = cr_in[10];
  assign n12925_o = cr_in[11];
  /* execute1.vhdl:719:39  */
  assign n12926_o = cr_in[12];
  assign n12927_o = cr_in[13];
  /* execute1.vhdl:719:29  */
  assign n12928_o = cr_in[14];
  assign n12929_o = cr_in[15];
  /* execute1.vhdl:719:29  */
  assign n12930_o = cr_in[16];
  /* execute1.vhdl:718:31  */
  assign n12931_o = cr_in[17];
  /* insn_helpers.vhdl:23:14  */
  assign n12932_o = cr_in[18];
  /* insn_helpers.vhdl:23:14  */
  assign n12933_o = cr_in[19];
  assign n12934_o = cr_in[20];
  /* insn_helpers.vhdl:23:14  */
  assign n12935_o = cr_in[21];
  assign n12936_o = cr_in[22];
  assign n12937_o = cr_in[23];
  /* insn_helpers.vhdl:27:14  */
  assign n12938_o = cr_in[24];
  /* insn_helpers.vhdl:27:14  */
  assign n12939_o = cr_in[25];
  assign n12940_o = cr_in[26];
  /* insn_helpers.vhdl:27:14  */
  assign n12941_o = cr_in[27];
  /* insn_helpers.vhdl:26:14  */
  assign n12942_o = cr_in[28];
  /* insn_helpers.vhdl:26:14  */
  assign n12943_o = cr_in[29];
  assign n12944_o = cr_in[30];
  /* insn_helpers.vhdl:26:14  */
  assign n12945_o = cr_in[31];
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12946_o = n11262_o[1:0];
  /* ppc_fx_insns.vhdl:827:43  */
  always @*
    case (n12946_o)
      2'b00: n12947_o = n12914_o;
      2'b01: n12947_o = n12915_o;
      2'b10: n12947_o = n12916_o;
      2'b11: n12947_o = n12917_o;
    endcase
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12948_o = n11262_o[1:0];
  /* ppc_fx_insns.vhdl:827:43  */
  always @*
    case (n12948_o)
      2'b00: n12949_o = n12918_o;
      2'b01: n12949_o = n12919_o;
      2'b10: n12949_o = n12920_o;
      2'b11: n12949_o = n12921_o;
    endcase
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12950_o = n11262_o[1:0];
  /* ppc_fx_insns.vhdl:827:43  */
  always @*
    case (n12950_o)
      2'b00: n12951_o = n12922_o;
      2'b01: n12951_o = n12923_o;
      2'b10: n12951_o = n12924_o;
      2'b11: n12951_o = n12925_o;
    endcase
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12952_o = n11262_o[1:0];
  /* ppc_fx_insns.vhdl:827:43  */
  always @*
    case (n12952_o)
      2'b00: n12953_o = n12926_o;
      2'b01: n12953_o = n12927_o;
      2'b10: n12953_o = n12928_o;
      2'b11: n12953_o = n12929_o;
    endcase
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12954_o = n11262_o[1:0];
  /* ppc_fx_insns.vhdl:827:43  */
  always @*
    case (n12954_o)
      2'b00: n12955_o = n12930_o;
      2'b01: n12955_o = n12931_o;
      2'b10: n12955_o = n12932_o;
      2'b11: n12955_o = n12933_o;
    endcase
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12956_o = n11262_o[1:0];
  /* ppc_fx_insns.vhdl:827:43  */
  always @*
    case (n12956_o)
      2'b00: n12957_o = n12934_o;
      2'b01: n12957_o = n12935_o;
      2'b10: n12957_o = n12936_o;
      2'b11: n12957_o = n12937_o;
    endcase
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12958_o = n11262_o[1:0];
  /* ppc_fx_insns.vhdl:827:43  */
  always @*
    case (n12958_o)
      2'b00: n12959_o = n12938_o;
      2'b01: n12959_o = n12939_o;
      2'b10: n12959_o = n12940_o;
      2'b11: n12959_o = n12941_o;
    endcase
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12960_o = n11262_o[1:0];
  /* ppc_fx_insns.vhdl:827:43  */
  always @*
    case (n12960_o)
      2'b00: n12961_o = n12942_o;
      2'b01: n12961_o = n12943_o;
      2'b10: n12961_o = n12944_o;
      2'b11: n12961_o = n12945_o;
    endcase
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12962_o = n11262_o[3:2];
  /* ppc_fx_insns.vhdl:827:43  */
  always @*
    case (n12962_o)
      2'b00: n12963_o = n12947_o;
      2'b01: n12963_o = n12949_o;
      2'b10: n12963_o = n12951_o;
      2'b11: n12963_o = n12953_o;
    endcase
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12964_o = n11262_o[3:2];
  /* ppc_fx_insns.vhdl:827:43  */
  always @*
    case (n12964_o)
      2'b00: n12965_o = n12955_o;
      2'b01: n12965_o = n12957_o;
      2'b10: n12965_o = n12959_o;
      2'b11: n12965_o = n12961_o;
    endcase
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12966_o = n11262_o[4];
  /* ppc_fx_insns.vhdl:827:43  */
  assign n12967_o = n12966_o ? n12965_o : n12963_o;
endmodule

module cr_file_0_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clk,
   input  d_in_read,
   input  w_in_write_cr_enable,
   input  [7:0] w_in_write_cr_mask,
   input  [31:0] w_in_write_cr_data,
   input  w_in_write_xerc_enable,
   input  [4:0] w_in_write_xerc_data,
   input  sim_dump,
   output [31:0] d_out_read_cr_data,
   output [4:0] d_out_read_xerc_data,
   output [12:0] log_out);
  wire [31:0] n9034_o;
  wire [4:0] n9035_o;
  wire [46:0] n9036_o;
  reg [31:0] crs;
  wire [31:0] crs_updated;
  reg [4:0] xerc;
  wire [4:0] xerc_updated;
  wire n9044_o;
  wire [3:0] n9045_o;
  wire [3:0] n9050_o;
  wire [3:0] n9051_o;
  wire n9053_o;
  wire [3:0] n9054_o;
  wire [3:0] n9059_o;
  wire [3:0] n9060_o;
  wire n9062_o;
  wire [3:0] n9063_o;
  wire [3:0] n9068_o;
  wire [3:0] n9069_o;
  wire n9071_o;
  wire [3:0] n9072_o;
  wire [3:0] n9077_o;
  wire [3:0] n9078_o;
  wire n9080_o;
  wire [3:0] n9081_o;
  wire [3:0] n9086_o;
  wire [3:0] n9087_o;
  wire n9089_o;
  wire [3:0] n9090_o;
  wire [3:0] n9095_o;
  wire [3:0] n9096_o;
  wire n9098_o;
  wire [3:0] n9099_o;
  wire [3:0] n9104_o;
  wire [3:0] n9105_o;
  wire [3:0] n9106_o;
  wire n9107_o;
  wire [3:0] n9108_o;
  wire [3:0] n9113_o;
  wire [31:0] n9114_o;
  wire n9115_o;
  wire [4:0] n9116_o;
  wire [4:0] n9117_o;
  wire n9122_o;
  wire n9124_o;
  wire [31:0] n9132_o;
  reg [31:0] n9133_q;
  wire [4:0] n9134_o;
  reg [4:0] n9135_q;
  wire [36:0] n9136_o;
  localparam [12:0] n9137_o = 13'bZ;
  assign d_out_read_cr_data = n9034_o;
  assign d_out_read_xerc_data = n9035_o;
  assign log_out = n9137_o;
  /* asic/register_file.vhdl:65:20  */
  assign n9034_o = n9136_o[31:0];
  /* asic/register_file.vhdl:30:9  */
  assign n9035_o = n9136_o[36:32];
  /* asic/register_file.vhdl:28:9  */
  assign n9036_o = {w_in_write_xerc_data, w_in_write_xerc_enable, w_in_write_cr_data, w_in_write_cr_mask, w_in_write_cr_enable};
  /* cr_file.vhdl:30:12  */
  always @*
    crs = n9133_q; // (isignal)
  initial
    crs = 32'b00000000000000000000000000000000;
  /* cr_file.vhdl:31:12  */
  assign crs_updated = n9114_o; // (signal)
  /* cr_file.vhdl:32:12  */
  always @*
    xerc = n9135_q; // (isignal)
  initial
    xerc = 5'b00000;
  /* cr_file.vhdl:33:12  */
  assign xerc_updated = n9117_o; // (signal)
  /* cr_file.vhdl:42:34  */
  assign n9044_o = n9036_o[1];
  /* cr_file.vhdl:45:59  */
  assign n9045_o = n9036_o[12:9];
  assign n9050_o = crs[3:0];
  /* cr_file.vhdl:42:13  */
  assign n9051_o = n9044_o ? n9045_o : n9050_o;
  /* cr_file.vhdl:42:34  */
  assign n9053_o = n9036_o[2];
  /* cr_file.vhdl:45:59  */
  assign n9054_o = n9036_o[16:13];
  /* common.vhdl:112:14  */
  assign n9059_o = crs[7:4];
  /* cr_file.vhdl:42:13  */
  assign n9060_o = n9053_o ? n9054_o : n9059_o;
  /* cr_file.vhdl:42:34  */
  assign n9062_o = n9036_o[3];
  /* cr_file.vhdl:45:59  */
  assign n9063_o = n9036_o[20:17];
  /* insn_helpers.vhdl:41:14  */
  assign n9068_o = crs[11:8];
  /* cr_file.vhdl:42:13  */
  assign n9069_o = n9062_o ? n9063_o : n9068_o;
  /* cr_file.vhdl:42:34  */
  assign n9071_o = n9036_o[4];
  /* cr_file.vhdl:45:59  */
  assign n9072_o = n9036_o[24:21];
  assign n9077_o = crs[15:12];
  /* cr_file.vhdl:42:13  */
  assign n9078_o = n9071_o ? n9072_o : n9077_o;
  /* cr_file.vhdl:42:34  */
  assign n9080_o = n9036_o[5];
  /* cr_file.vhdl:45:59  */
  assign n9081_o = n9036_o[28:25];
  /* insn_helpers.vhdl:6:14  */
  assign n9086_o = crs[19:16];
  /* cr_file.vhdl:42:13  */
  assign n9087_o = n9080_o ? n9081_o : n9086_o;
  /* cr_file.vhdl:42:34  */
  assign n9089_o = n9036_o[6];
  /* cr_file.vhdl:45:59  */
  assign n9090_o = n9036_o[32:29];
  /* insn_helpers.vhdl:44:14  */
  assign n9095_o = crs[23:20];
  /* cr_file.vhdl:42:13  */
  assign n9096_o = n9089_o ? n9090_o : n9095_o;
  /* cr_file.vhdl:42:34  */
  assign n9098_o = n9036_o[7];
  /* cr_file.vhdl:45:59  */
  assign n9099_o = n9036_o[36:33];
  /* insn_helpers.vhdl:41:14  */
  assign n9104_o = crs[27:24];
  /* cr_file.vhdl:42:13  */
  assign n9105_o = n9098_o ? n9099_o : n9104_o;
  /* insn_helpers.vhdl:41:14  */
  assign n9106_o = crs[31:28];
  /* cr_file.vhdl:42:34  */
  assign n9107_o = n9036_o[8];
  /* cr_file.vhdl:45:59  */
  assign n9108_o = n9036_o[40:37];
  /* cr_file.vhdl:42:13  */
  assign n9113_o = n9107_o ? n9108_o : n9106_o;
  /* insn_helpers.vhdl:9:14  */
  assign n9114_o = {n9113_o, n9105_o, n9096_o, n9087_o, n9078_o, n9069_o, n9060_o, n9051_o};
  /* cr_file.vhdl:51:17  */
  assign n9115_o = n9036_o[41];
  /* cr_file.vhdl:52:34  */
  assign n9116_o = n9036_o[46:42];
  /* cr_file.vhdl:51:9  */
  assign n9117_o = n9115_o ? n9116_o : xerc;
  /* cr_file.vhdl:63:21  */
  assign n9122_o = n9036_o[0];
  /* cr_file.vhdl:67:21  */
  assign n9124_o = n9036_o[41];
  /* cr_file.vhdl:62:9  */
  assign n9132_o = n9122_o ? crs_updated : crs;
  /* cr_file.vhdl:62:9  */
  always @(posedge clk)
    n9133_q <= n9132_o;
  initial
    n9133_q = 32'b00000000000000000000000000000000;
  /* cr_file.vhdl:62:9  */
  assign n9134_o = n9124_o ? xerc_updated : xerc;
  /* cr_file.vhdl:62:9  */
  always @(posedge clk)
    n9135_q <= n9134_o;
  initial
    n9135_q = 5'b00000;
  /* cr_file.vhdl:62:9  */
  assign n9136_o = {xerc_updated, crs_updated};
endmodule

module register_file_0_3f29546453678b855931c174a97d6c0894b8f546
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  clk,
   input  d_in_read1_enable,
   input  [6:0] d_in_read1_reg,
   input  d_in_read2_enable,
   input  [6:0] d_in_read2_reg,
   input  d_in_read3_enable,
   input  [6:0] d_in_read3_reg,
   input  [6:0] w_in_write_reg,
   input  [63:0] w_in_write_data,
   input  w_in_write_enable,
   input  dbg_gpr_req,
   input  [6:0] dbg_gpr_addr,
   input  sim_dump,
   output [63:0] d_out_read1_data,
   output [63:0] d_out_read2_data,
   output [63:0] d_out_read3_data,
   output dbg_gpr_ack,
   output [63:0] dbg_gpr_data,
   output sim_dump_done,
   output [71:0] log_out);
  wire [23:0] n8985_o;
  wire [63:0] n8987_o;
  wire [63:0] n8988_o;
  wire [63:0] n8989_o;
  wire [71:0] n8990_o;
  wire [63:0] d1;
  wire [63:0] d2;
  wire [63:0] d3;
  wire [63:0] register_file_0_D1;
  wire [63:0] register_file_0_D2;
  wire [63:0] register_file_0_D3;
  wire [6:0] n8995_o;
  wire [6:0] n8996_o;
  wire [6:0] n8997_o;
  wire n9001_o;
  wire [6:0] n9002_o;
  wire [63:0] n9003_o;
  wire n9009_o;
  wire [6:0] n9010_o;
  wire [6:0] n9011_o;
  wire n9012_o;
  wire [63:0] n9013_o;
  wire [63:0] n9014_o;
  wire [6:0] n9015_o;
  wire [6:0] n9016_o;
  wire n9017_o;
  wire [63:0] n9018_o;
  wire [63:0] n9019_o;
  wire [6:0] n9020_o;
  wire [6:0] n9021_o;
  wire n9022_o;
  wire [63:0] n9023_o;
  wire [63:0] n9024_o;
  wire [191:0] n9025_o;
  wire [191:0] n9026_o;
  wire [191:0] n9027_o;
  localparam n9029_o = 1'bZ;
  localparam [63:0] n9030_o = 64'bZ;
  localparam n9031_o = 1'bZ;
  localparam [71:0] n9032_o = 72'bZ;
  assign d_out_read1_data = n8987_o;
  assign d_out_read2_data = n8988_o;
  assign d_out_read3_data = n8989_o;
  assign dbg_gpr_ack = n9029_o;
  assign dbg_gpr_data = n9030_o;
  assign sim_dump_done = n9031_o;
  assign log_out = n9032_o;
  /* decode2.vhdl:345:30  */
  assign n8985_o = {d_in_read3_reg, d_in_read3_enable, d_in_read2_reg, d_in_read2_enable, d_in_read1_reg, d_in_read1_enable};
  /* decode2.vhdl:343:29  */
  assign n8987_o = n9027_o[63:0];
  /* decode2.vhdl:342:29  */
  assign n8988_o = n9027_o[127:64];
  /* decode2.vhdl:341:29  */
  assign n8989_o = n9027_o[191:128];
  /* decode2.vhdl:339:28  */
  assign n8990_o = {w_in_write_enable, w_in_write_data, w_in_write_reg};
  /* asic/register_file.vhdl:52:12  */
  assign d1 = register_file_0_D1; // (signal)
  /* asic/register_file.vhdl:53:12  */
  assign d2 = register_file_0_D2; // (signal)
  /* asic/register_file.vhdl:54:12  */
  assign d3 = register_file_0_D3; // (signal)
  /* asic/register_file.vhdl:57:5  */
  Microwatt_FP_DFFRFile register_file_0 (
`ifdef USE_POWER_PINS
    .VPWR(vccd1),
    .VGND(vssd1),
`endif
    .CLK(clk),
    .R1(n8995_o),
    .R2(n8996_o),
    .R3(n8997_o),
    .WE(n9001_o),
    .RW(n9002_o),
    .DW(n9003_o),
    .D1(register_file_0_D1),
    .D2(register_file_0_D2),
    .D3(register_file_0_D3));
  /* asic/register_file.vhdl:61:25  */
  assign n8995_o = n8985_o[7:1];
  /* asic/register_file.vhdl:62:25  */
  assign n8996_o = n8985_o[15:9];
  /* asic/register_file.vhdl:63:25  */
  assign n8997_o = n8985_o[23:17];
  /* asic/register_file.vhdl:69:25  */
  assign n9001_o = n8990_o[71];
  /* asic/register_file.vhdl:70:25  */
  assign n9002_o = n8990_o[6:0];
  /* asic/register_file.vhdl:71:25  */
  assign n9003_o = n8990_o[70:7];
  /* asic/register_file.vhdl:90:17  */
  assign n9009_o = n8990_o[71];
  /* asic/register_file.vhdl:91:21  */
  assign n9010_o = n8985_o[7:1];
  /* asic/register_file.vhdl:91:38  */
  assign n9011_o = n8990_o[6:0];
  /* asic/register_file.vhdl:91:31  */
  assign n9012_o = n9010_o == n9011_o;
  /* asic/register_file.vhdl:92:42  */
  assign n9013_o = n8990_o[70:7];
  /* asic/register_file.vhdl:91:13  */
  assign n9014_o = n9012_o ? n9013_o : d1;
  /* asic/register_file.vhdl:94:21  */
  assign n9015_o = n8985_o[15:9];
  /* asic/register_file.vhdl:94:38  */
  assign n9016_o = n8990_o[6:0];
  /* asic/register_file.vhdl:94:31  */
  assign n9017_o = n9015_o == n9016_o;
  /* asic/register_file.vhdl:95:42  */
  assign n9018_o = n8990_o[70:7];
  /* asic/register_file.vhdl:94:13  */
  assign n9019_o = n9017_o ? n9018_o : d2;
  /* asic/register_file.vhdl:97:21  */
  assign n9020_o = n8985_o[23:17];
  /* asic/register_file.vhdl:97:38  */
  assign n9021_o = n8990_o[6:0];
  /* asic/register_file.vhdl:97:31  */
  assign n9022_o = n9020_o == n9021_o;
  /* asic/register_file.vhdl:98:42  */
  assign n9023_o = n8990_o[70:7];
  /* asic/register_file.vhdl:97:13  */
  assign n9024_o = n9022_o ? n9023_o : d3;
  assign n9025_o = {n9024_o, n9019_o, n9014_o};
  /* insn_helpers.vhdl:19:14  */
  assign n9026_o = {d3, d2, d1};
  /* asic/register_file.vhdl:90:9  */
  assign n9027_o = n9009_o ? n9025_o : n9026_o;
endmodule

module decode2_0_9159cb8bcee7fcb95582f140960cdae72788d326
  (input  clk,
   input  rst,
   input  [1:0] complete_in_tag,
   input  complete_in_valid,
   input  busy_in,
   input  flush_in,
   input  d_in_valid,
   input  d_in_stop_mark,
   input  [63:0] d_in_nia,
   input  [31:0] d_in_insn,
   input  [6:0] d_in_ispr1,
   input  [6:0] d_in_ispr2,
   input  [6:0] d_in_ispro,
   input  [43:0] d_in_decode,
   input  d_in_br_pred,
   input  d_in_big_endian,
   input  [63:0] r_in_read1_data,
   input  [63:0] r_in_read2_data,
   input  [63:0] r_in_read3_data,
   input  [31:0] c_in_read_cr_data,
   input  [4:0] c_in_read_xerc_data,
   input  [2:0] execute_bypass_tag,
   input  [63:0] execute_bypass_data,
   input  [2:0] execute_cr_bypass_tag,
   input  [31:0] execute_cr_bypass_data,
   output stall_out,
   output stopped_out,
   output e_out_valid,
   output [1:0] e_out_unit,
   output e_out_fac,
   output [5:0] e_out_insn_type,
   output [63:0] e_out_nia,
   output [2:0] e_out_instr_tag,
   output [6:0] e_out_write_reg,
   output e_out_write_reg_enable,
   output [6:0] e_out_read_reg1,
   output [6:0] e_out_read_reg2,
   output [63:0] e_out_read_data1,
   output [63:0] e_out_read_data2,
   output [63:0] e_out_read_data3,
   output [31:0] e_out_cr,
   output [4:0] e_out_xerc,
   output e_out_lr,
   output e_out_br_abs,
   output e_out_rc,
   output e_out_oe,
   output e_out_invert_a,
   output e_out_addm1,
   output e_out_invert_out,
   output [1:0] e_out_input_carry,
   output e_out_output_carry,
   output e_out_input_cr,
   output e_out_output_cr,
   output e_out_output_xer,
   output e_out_is_32bit,
   output e_out_is_signed,
   output [31:0] e_out_insn,
   output [3:0] e_out_data_len,
   output e_out_byte_reverse,
   output e_out_sign_extend,
   output e_out_update,
   output e_out_reserve,
   output e_out_br_pred,
   output [2:0] e_out_result_sel,
   output [2:0] e_out_sub_select,
   output e_out_repeat,
   output e_out_second,
   output r_out_read1_enable,
   output [6:0] r_out_read1_reg,
   output r_out_read2_enable,
   output [6:0] r_out_read2_reg,
   output r_out_read3_enable,
   output [6:0] r_out_read3_reg,
   output c_out_read,
   output [9:0] log_out);
  wire [2:0] n8029_o;
  wire [164:0] n8032_o;
  wire n8034_o;
  wire [1:0] n8035_o;
  wire n8036_o;
  wire [5:0] n8037_o;
  wire [63:0] n8038_o;
  wire [2:0] n8039_o;
  wire [6:0] n8040_o;
  wire n8041_o;
  wire [6:0] n8042_o;
  wire [6:0] n8043_o;
  wire [63:0] n8044_o;
  wire [63:0] n8045_o;
  wire [63:0] n8046_o;
  wire [31:0] n8047_o;
  wire [4:0] n8048_o;
  wire n8049_o;
  wire n8050_o;
  wire n8051_o;
  wire n8052_o;
  wire n8053_o;
  wire n8054_o;
  wire n8055_o;
  wire [1:0] n8056_o;
  wire n8057_o;
  wire n8058_o;
  wire n8059_o;
  wire n8060_o;
  wire n8061_o;
  wire n8062_o;
  wire [31:0] n8063_o;
  wire [3:0] n8064_o;
  wire n8065_o;
  wire n8066_o;
  wire n8067_o;
  wire n8068_o;
  wire n8069_o;
  wire [2:0] n8070_o;
  wire [2:0] n8071_o;
  wire n8072_o;
  wire n8073_o;
  wire [191:0] n8074_o;
  wire n8076_o;
  wire [6:0] n8077_o;
  wire n8078_o;
  wire [6:0] n8079_o;
  wire n8080_o;
  wire [6:0] n8081_o;
  wire [36:0] n8082_o;
  wire n8084_o;
  wire [66:0] n8085_o;
  wire [34:0] n8086_o;
  wire [392:0] r;
  wire [392:0] rin;
  wire deferred;
  wire control_valid_in;
  wire control_valid_out;
  wire control_stall_out;
  wire control_sgl_pipe;
  wire gpr_write_valid;
  wire [6:0] gpr_write;
  wire gpr_a_read_valid;
  wire [6:0] gpr_a_read;
  wire gpr_a_bypass;
  wire gpr_b_read_valid;
  wire [6:0] gpr_b_read;
  wire gpr_b_bypass;
  wire gpr_c_read_valid;
  wire [6:0] gpr_c_read;
  wire gpr_c_bypass;
  wire cr_read_valid;
  wire cr_write_valid;
  wire cr_bypass;
  wire [2:0] instr_tag;
  wire control_0_valid_out;
  wire control_0_stall_out;
  wire control_0_stopped_out;
  wire control_0_gpr_bypass_a;
  wire control_0_gpr_bypass_b;
  wire control_0_gpr_bypass_c;
  wire control_0_cr_bypass;
  wire [1:0] control_0_instr_tag_out_tag;
  wire control_0_instr_tag_out_valid;
  wire [1:0] n8088_o;
  wire n8089_o;
  wire n8090_o;
  wire n8091_o;
  wire [2:0] n8092_o;
  wire [1:0] n8093_o;
  wire n8094_o;
  wire [2:0] n8095_o;
  wire [1:0] n8096_o;
  wire n8097_o;
  wire [2:0] n8105_o;
  wire [391:0] n8107_o;
  wire n8108_o;
  wire n8109_o;
  wire n8112_o;
  wire n8113_o;
  wire n8114_o;
  wire [43:0] n8120_o;
  wire n8121_o;
  localparam [391:0] n8132_o = 392'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire n8133_o;
  wire [43:0] n8134_o;
  wire n8135_o;
  wire [43:0] n8138_o;
  wire n8139_o;
  wire [50:0] n8140_o;
  wire [43:0] n8141_o;
  wire [5:0] n8142_o;
  wire [5:0] n8143_o;
  wire n8145_o;
  wire [31:0] n8147_o;
  wire n8152_o;
  wire n8153_o;
  wire n8156_o;
  wire n8157_o;
  wire n8158_o;
  wire n8160_o;
  wire n8162_o;
  wire n8163_o;
  wire n8165_o;
  wire n8166_o;
  wire n8168_o;
  wire n8169_o;
  wire [31:0] n8171_o;
  wire [4:0] n8176_o;
  wire [4:0] n8177_o;
  wire [9:0] n8178_o;
  wire [31:0] n8180_o;
  wire n8182_o;
  wire n8184_o;
  wire n8186_o;
  wire [1:0] n8187_o;
  wire n8188_o;
  reg n8189_o;
  reg n8190_o;
  wire [6:0] n8191_o;
  wire [43:0] n8194_o;
  wire [2:0] n8195_o;
  wire [31:0] n8196_o;
  wire [63:0] n8197_o;
  wire [6:0] n8198_o;
  wire [63:0] n8199_o;
  wire n8205_o;
  wire n8207_o;
  wire [4:0] n8213_o;
  wire n8215_o;
  wire n8216_o;
  wire n8217_o;
  wire [4:0] n8224_o;
  wire [6:0] n8230_o;
  wire [71:0] n8232_o;
  wire n8234_o;
  wire n8240_o;
  wire [71:0] n8241_o;
  wire n8243_o;
  wire [71:0] n8246_o;
  wire n8248_o;
  wire n8250_o;
  wire [4:0] n8257_o;
  wire [6:0] n8263_o;
  wire [71:0] n8265_o;
  wire [71:0] n8267_o;
  wire [71:0] n8268_o;
  wire [71:0] n8269_o;
  wire [71:0] n8270_o;
  wire [43:0] n8272_o;
  wire [3:0] n8273_o;
  wire [31:0] n8274_o;
  wire [63:0] n8275_o;
  wire [6:0] n8276_o;
  wire [4:0] n8288_o;
  wire [6:0] n8294_o;
  wire [71:0] n8296_o;
  wire n8298_o;
  wire [4:0] n8305_o;
  wire [6:0] n8311_o;
  wire [71:0] n8313_o;
  wire n8315_o;
  wire [15:0] n8321_o;
  wire [63:0] n8322_o;
  wire [71:0] n8325_o;
  wire n8327_o;
  wire [15:0] n8333_o;
  wire [63:0] n8334_o;
  wire [71:0] n8337_o;
  wire n8339_o;
  wire [15:0] n8345_o;
  wire [31:0] n8347_o;
  wire [63:0] n8348_o;
  wire [71:0] n8351_o;
  wire n8353_o;
  wire [15:0] n8359_o;
  wire [31:0] n8361_o;
  wire [63:0] n8362_o;
  wire [71:0] n8365_o;
  wire n8367_o;
  wire [23:0] n8373_o;
  wire [25:0] n8375_o;
  wire [63:0] n8376_o;
  wire [71:0] n8379_o;
  wire n8381_o;
  wire [13:0] n8387_o;
  wire [15:0] n8389_o;
  wire [63:0] n8390_o;
  wire [71:0] n8393_o;
  wire n8395_o;
  wire [13:0] n8401_o;
  wire [15:0] n8403_o;
  wire [63:0] n8404_o;
  wire [71:0] n8407_o;
  wire n8409_o;
  wire [11:0] n8415_o;
  wire [15:0] n8417_o;
  wire [63:0] n8418_o;
  wire [71:0] n8421_o;
  wire n8423_o;
  wire [9:0] n8429_o;
  wire [4:0] n8430_o;
  wire [14:0] n8431_o;
  wire n8432_o;
  wire [15:0] n8433_o;
  wire [31:0] n8435_o;
  wire [63:0] n8436_o;
  wire [71:0] n8439_o;
  wire n8441_o;
  wire n8443_o;
  wire n8444_o;
  wire [58:0] n8446_o;
  wire [4:0] n8447_o;
  wire [63:0] n8448_o;
  wire [71:0] n8451_o;
  wire n8453_o;
  wire [4:0] n8454_o;
  wire [63:0] n8456_o;
  wire [71:0] n8459_o;
  wire n8461_o;
  wire n8467_o;
  wire [71:0] n8468_o;
  wire n8470_o;
  wire n8472_o;
  wire [15:0] n8473_o;
  reg [71:0] n8477_o;
  wire [43:0] n8480_o;
  wire [2:0] n8481_o;
  wire [31:0] n8482_o;
  wire [63:0] n8483_o;
  wire [4:0] n8494_o;
  wire [6:0] n8500_o;
  wire [71:0] n8502_o;
  wire n8504_o;
  wire [4:0] n8511_o;
  wire [6:0] n8517_o;
  wire [71:0] n8519_o;
  wire n8521_o;
  wire [4:0] n8528_o;
  wire [6:0] n8534_o;
  wire [71:0] n8536_o;
  wire n8538_o;
  wire [4:0] n8545_o;
  wire [6:0] n8551_o;
  wire [71:0] n8553_o;
  wire n8555_o;
  wire n8558_o;
  wire [4:0] n8559_o;
  reg [71:0] n8561_o;
  wire [43:0] n8563_o;
  wire [2:0] n8564_o;
  wire [31:0] n8565_o;
  wire [6:0] n8566_o;
  wire [4:0] n8577_o;
  wire [6:0] n8583_o;
  wire [7:0] n8585_o;
  wire n8587_o;
  wire [4:0] n8594_o;
  wire [6:0] n8600_o;
  wire [7:0] n8602_o;
  wire n8604_o;
  wire [4:0] n8611_o;
  wire [6:0] n8617_o;
  wire [7:0] n8619_o;
  wire n8621_o;
  wire n8627_o;
  wire [7:0] n8628_o;
  wire n8630_o;
  wire n8633_o;
  wire [4:0] n8634_o;
  reg [7:0] n8636_o;
  wire [43:0] n8637_o;
  wire n8638_o;
  wire [31:0] n8640_o;
  wire n8645_o;
  wire [31:0] n8647_o;
  wire n8652_o;
  wire n8653_o;
  wire n8654_o;
  wire [1:0] n8655_o;
  wire [1:0] n8656_o;
  wire [1:0] n8657_o;
  wire n8658_o;
  wire [327:0] n8659_o;
  wire [43:0] n8660_o;
  wire [5:0] n8661_o;
  wire [43:0] n8662_o;
  wire [1:0] n8663_o;
  wire n8665_o;
  wire n8667_o;
  wire [43:0] n8668_o;
  wire [1:0] n8669_o;
  wire n8670_o;
  wire n8671_o;
  wire n8672_o;
  wire n8674_o;
  wire n8675_o;
  wire n8677_o;
  wire n8678_o;
  wire n8679_o;
  wire n8680_o;
  wire n8682_o;
  wire n8683_o;
  wire n8685_o;
  wire n8686_o;
  wire [6:0] n8687_o;
  wire [6:0] n8688_o;
  wire [6:0] n8689_o;
  wire n8691_o;
  wire [2:0] n8692_o;
  wire n8693_o;
  reg n8694_o;
  wire n8695_o;
  wire n8696_o;
  reg n8697_o;
  wire [5:0] n8698_o;
  wire [5:0] n8699_o;
  reg [5:0] n8700_o;
  wire [392:0] n8701_o;
  wire [391:0] n8702_o;
  wire n8703_o;
  wire n8704_o;
  wire n8705_o;
  wire n8707_o;
  wire n8708_o;
  wire n8709_o;
  wire [1:0] n8710_o;
  wire [1:0] n8711_o;
  wire [1:0] n8712_o;
  wire n8713_o;
  wire n8714_o;
  wire [1:0] n8715_o;
  wire [1:0] n8716_o;
  wire n8718_o;
  wire n8719_o;
  wire [69:0] n8720_o;
  wire n8721_o;
  wire [6:0] n8722_o;
  wire n8723_o;
  wire n8724_o;
  wire [5:0] n8725_o;
  wire [5:0] n8726_o;
  wire [5:0] n8727_o;
  wire n8729_o;
  wire n8730_o;
  wire n8731_o;
  wire n8732_o;
  wire [6:0] n8733_o;
  wire n8734_o;
  wire n8735_o;
  wire n8736_o;
  wire [6:0] n8737_o;
  wire [71:0] n8738_o;
  wire n8739_o;
  wire n8740_o;
  wire n8741_o;
  wire [71:0] n8742_o;
  wire [6:0] n8743_o;
  wire [43:0] n8744_o;
  wire [2:0] n8745_o;
  wire n8747_o;
  wire n8749_o;
  wire n8751_o;
  wire n8753_o;
  wire n8755_o;
  wire [4:0] n8756_o;
  reg [3:0] n8763_o;
  wire [63:0] n8764_o;
  wire [43:0] n8767_o;
  wire [1:0] n8768_o;
  wire n8770_o;
  wire [43:0] n8771_o;
  wire n8772_o;
  wire [6:0] n8775_o;
  wire [6:0] n8778_o;
  wire [7:0] n8780_o;
  wire [6:0] n8781_o;
  wire [7:0] n8783_o;
  wire n8784_o;
  wire [43:0] n8786_o;
  wire [1:0] n8787_o;
  wire [31:0] n8788_o;
  wire n8798_o;
  wire n8800_o;
  wire n8803_o;
  wire n8806_o;
  wire [2:0] n8807_o;
  reg n8809_o;
  wire [4:0] n8810_o;
  wire [43:0] n8812_o;
  wire n8813_o;
  wire [43:0] n8817_o;
  wire n8818_o;
  wire [43:0] n8820_o;
  wire [1:0] n8821_o;
  wire [43:0] n8823_o;
  wire n8824_o;
  wire n8825_o;
  wire [43:0] n8826_o;
  wire n8827_o;
  wire [43:0] n8829_o;
  wire n8830_o;
  wire [31:0] n8832_o;
  wire [43:0] n8835_o;
  wire n8836_o;
  wire [43:0] n8838_o;
  wire n8839_o;
  wire [43:0] n8841_o;
  wire n8842_o;
  wire [43:0] n8844_o;
  wire n8845_o;
  wire n8847_o;
  wire [5:0] n8850_o;
  wire [5:0] n8856_o;
  wire n8861_o;
  wire n8863_o;
  wire n8864_o;
  wire n8865_o;
  wire n8866_o;
  wire n8867_o;
  wire n8868_o;
  wire n8869_o;
  wire [43:0] n8870_o;
  wire [5:0] n8871_o;
  wire n8873_o;
  wire n8874_o;
  wire n8875_o;
  wire n8876_o;
  wire n8877_o;
  wire n8878_o;
  wire n8881_o;
  wire [2:0] n8882_o;
  wire n8883_o;
  wire n8884_o;
  wire [63:0] n8885_o;
  wire n8887_o;
  wire [63:0] n8888_o;
  reg [63:0] n8889_o;
  wire [63:0] n8891_o;
  wire n8893_o;
  wire [63:0] n8894_o;
  reg [63:0] n8895_o;
  wire [63:0] n8897_o;
  wire n8899_o;
  wire [71:0] n8900_o;
  wire [63:0] n8901_o;
  reg [63:0] n8902_o;
  wire [31:0] n8904_o;
  wire [31:0] n8905_o;
  wire [31:0] n8906_o;
  wire n8907_o;
  wire [43:0] n8908_o;
  wire n8909_o;
  wire [392:0] n8910_o;
  wire [391:0] n8911_o;
  wire n8912_o;
  wire [7:0] n8913_o;
  wire [6:0] n8914_o;
  wire n8915_o;
  wire [6:0] n8916_o;
  wire n8917_o;
  wire [6:0] n8918_o;
  wire [71:0] n8919_o;
  wire n8920_o;
  wire [71:0] n8921_o;
  wire [6:0] n8922_o;
  wire [43:0] n8923_o;
  wire n8924_o;
  wire [43:0] n8926_o;
  wire [1:0] n8927_o;
  wire [31:0] n8928_o;
  wire n8938_o;
  wire n8940_o;
  wire n8943_o;
  wire n8946_o;
  wire [2:0] n8947_o;
  reg n8949_o;
  wire n8950_o;
  wire [43:0] n8951_o;
  wire n8952_o;
  wire n8953_o;
  wire [392:0] n8954_o;
  wire [391:0] n8955_o;
  wire n8956_o;
  wire n8957_o;
  wire n8958_o;
  wire n8959_o;
  wire n8960_o;
  wire [392:0] n8961_o;
  wire n8962_o;
  wire n8963_o;
  wire n8964_o;
  wire [392:0] n8967_o;
  wire [392:0] n8968_o;
  wire [392:0] n8969_o;
  wire [391:0] n8970_o;
  wire [392:0] n8977_o;
  reg [392:0] n8978_q;
  wire [23:0] n8979_o;
  localparam [9:0] n8980_o = 10'bZ;
  wire [2:0] n8982_data; // mem_rd
  wire [2:0] n8984_data; // mem_rd
  assign stall_out = n8963_o;
  assign stopped_out = control_0_stopped_out;
  assign e_out_valid = n8034_o;
  assign e_out_unit = n8035_o;
  assign e_out_fac = n8036_o;
  assign e_out_insn_type = n8037_o;
  assign e_out_nia = n8038_o;
  assign e_out_instr_tag = n8039_o;
  assign e_out_write_reg = n8040_o;
  assign e_out_write_reg_enable = n8041_o;
  assign e_out_read_reg1 = n8042_o;
  assign e_out_read_reg2 = n8043_o;
  assign e_out_read_data1 = n8044_o;
  assign e_out_read_data2 = n8045_o;
  assign e_out_read_data3 = n8046_o;
  assign e_out_cr = n8047_o;
  assign e_out_xerc = n8048_o;
  assign e_out_lr = n8049_o;
  assign e_out_br_abs = n8050_o;
  assign e_out_rc = n8051_o;
  assign e_out_oe = n8052_o;
  assign e_out_invert_a = n8053_o;
  assign e_out_addm1 = n8054_o;
  assign e_out_invert_out = n8055_o;
  assign e_out_input_carry = n8056_o;
  assign e_out_output_carry = n8057_o;
  assign e_out_input_cr = n8058_o;
  assign e_out_output_cr = n8059_o;
  assign e_out_output_xer = n8060_o;
  assign e_out_is_32bit = n8061_o;
  assign e_out_is_signed = n8062_o;
  assign e_out_insn = n8063_o;
  assign e_out_data_len = n8064_o;
  assign e_out_byte_reverse = n8065_o;
  assign e_out_sign_extend = n8066_o;
  assign e_out_update = n8067_o;
  assign e_out_reserve = n8068_o;
  assign e_out_br_pred = n8069_o;
  assign e_out_result_sel = n8070_o;
  assign e_out_sub_select = n8071_o;
  assign e_out_repeat = n8072_o;
  assign e_out_second = n8073_o;
  assign r_out_read1_enable = n8076_o;
  assign r_out_read1_reg = n8077_o;
  assign r_out_read2_enable = n8078_o;
  assign r_out_read2_reg = n8079_o;
  assign r_out_read3_enable = n8080_o;
  assign r_out_read3_reg = n8081_o;
  assign c_out_read = n8084_o;
  assign log_out = n8980_o;
  /* decode1.vhdl:26:9  */
  assign n8029_o = {complete_in_valid, complete_in_tag};
  /* decode1.vhdl:21:9  */
  assign n8032_o = {d_in_big_endian, d_in_br_pred, d_in_decode, d_in_ispro, d_in_ispr2, d_in_ispr1, d_in_insn, d_in_nia, d_in_stop_mark, d_in_valid};
  /* decode1.vhdl:525:9  */
  assign n8034_o = n8970_o[0];
  assign n8035_o = n8970_o[2:1];
  assign n8036_o = n8970_o[3];
  assign n8037_o = n8970_o[9:4];
  assign n8038_o = n8970_o[73:10];
  assign n8039_o = n8970_o[76:74];
  /* decode1.vhdl:757:9  */
  assign n8040_o = n8970_o[83:77];
  assign n8041_o = n8970_o[84];
  assign n8042_o = n8970_o[91:85];
  assign n8043_o = n8970_o[98:92];
  /* decode1.vhdl:589:9  */
  assign n8044_o = n8970_o[162:99];
  /* decode1.vhdl:589:9  */
  assign n8045_o = n8970_o[226:163];
  /* decode1.vhdl:589:9  */
  assign n8046_o = n8970_o[290:227];
  assign n8047_o = n8970_o[322:291];
  assign n8048_o = n8970_o[327:323];
  assign n8049_o = n8970_o[328];
  assign n8050_o = n8970_o[329];
  assign n8051_o = n8970_o[330];
  assign n8052_o = n8970_o[331];
  /* decode1.vhdl:716:53  */
  assign n8053_o = n8970_o[332];
  /* decode1.vhdl:714:53  */
  assign n8054_o = n8970_o[333];
  /* decode1.vhdl:708:44  */
  assign n8055_o = n8970_o[334];
  /* decode1.vhdl:701:48  */
  assign n8056_o = n8970_o[336:335];
  /* decode1.vhdl:696:44  */
  assign n8057_o = n8970_o[337];
  /* decode1.vhdl:687:44  */
  assign n8058_o = n8970_o[338];
  /* decode1.vhdl:650:44  */
  assign n8059_o = n8970_o[339];
  /* decode1.vhdl:648:51  */
  assign n8060_o = n8970_o[340];
  /* common.vhdl:112:14  */
  assign n8061_o = n8970_o[341];
  /* common.vhdl:112:14  */
  assign n8062_o = n8970_o[342];
  assign n8063_o = n8970_o[374:343];
  /* common.vhdl:112:14  */
  assign n8064_o = n8970_o[378:375];
  /* common.vhdl:751:8  */
  assign n8065_o = n8970_o[379];
  assign n8066_o = n8970_o[380];
  /* common.vhdl:751:8  */
  assign n8067_o = n8970_o[381];
  assign n8068_o = n8970_o[382];
  assign n8069_o = n8970_o[383];
  /* common.vhdl:750:45  */
  assign n8070_o = n8970_o[386:384];
  assign n8071_o = n8970_o[389:387];
  assign n8072_o = n8970_o[390];
  /* common.vhdl:717:8  */
  assign n8073_o = n8970_o[391];
  assign n8074_o = {r_in_read3_data, r_in_read2_data, r_in_read1_data};
  assign n8076_o = n8979_o[0];
  /* common.vhdl:715:17  */
  assign n8077_o = n8979_o[7:1];
  assign n8078_o = n8979_o[8];
  /* common.vhdl:711:17  */
  assign n8079_o = n8979_o[15:9];
  assign n8080_o = n8979_o[16];
  /* common.vhdl:106:14  */
  assign n8081_o = n8979_o[23:17];
  /* common.vhdl:106:14  */
  assign n8082_o = {c_in_read_xerc_data, c_in_read_cr_data};
  /* common.vhdl:751:8  */
  assign n8084_o = n8121_o;
  assign n8085_o = {execute_bypass_data, execute_bypass_tag};
  /* common.vhdl:751:8  */
  assign n8086_o = {execute_cr_bypass_data, execute_cr_bypass_tag};
  /* decode2.vhdl:53:12  */
  assign r = n8978_q; // (signal)
  /* decode2.vhdl:53:15  */
  assign rin = n8969_o; // (signal)
  /* decode2.vhdl:55:12  */
  assign deferred = n8109_o; // (signal)
  /* decode2.vhdl:274:12  */
  assign control_valid_in = n8907_o; // (signal)
  /* decode2.vhdl:275:12  */
  assign control_valid_out = control_0_valid_out; // (signal)
  /* decode2.vhdl:276:12  */
  assign control_stall_out = control_0_stall_out; // (signal)
  /* decode2.vhdl:277:12  */
  assign control_sgl_pipe = n8909_o; // (signal)
  /* decode2.vhdl:279:12  */
  assign gpr_write_valid = n8912_o; // (signal)
  /* decode2.vhdl:280:12  */
  assign gpr_write = n8914_o; // (signal)
  /* decode2.vhdl:282:12  */
  assign gpr_a_read_valid = n8915_o; // (signal)
  /* decode2.vhdl:283:12  */
  assign gpr_a_read = n8916_o; // (signal)
  /* decode2.vhdl:284:12  */
  assign gpr_a_bypass = control_0_gpr_bypass_a; // (signal)
  /* decode2.vhdl:286:12  */
  assign gpr_b_read_valid = n8917_o; // (signal)
  /* decode2.vhdl:287:12  */
  assign gpr_b_read = n8918_o; // (signal)
  /* decode2.vhdl:288:12  */
  assign gpr_b_bypass = control_0_gpr_bypass_b; // (signal)
  /* decode2.vhdl:290:12  */
  assign gpr_c_read_valid = n8920_o; // (signal)
  /* decode2.vhdl:291:12  */
  assign gpr_c_read = n8922_o; // (signal)
  /* decode2.vhdl:292:12  */
  assign gpr_c_bypass = control_0_gpr_bypass_c; // (signal)
  /* decode2.vhdl:294:12  */
  assign cr_read_valid = n8953_o; // (signal)
  /* decode2.vhdl:295:12  */
  assign cr_write_valid = n8950_o; // (signal)
  /* decode2.vhdl:296:12  */
  assign cr_bypass = control_0_cr_bypass; // (signal)
  /* decode2.vhdl:298:12  */
  assign instr_tag = n8105_o; // (signal)
  /* decode2.vhdl:301:5  */
  control_3_bf8b4530d8d246dd74ac53a13471bba17941dff7 control_0 (
    .clk(clk),
    .rst(rst),
    .complete_in_tag(n8088_o),
    .complete_in_valid(n8089_o),
    .valid_in(control_valid_in),
    .repeated(n8090_o),
    .flush_in(flush_in),
    .busy_in(busy_in),
    .deferred(deferred),
    .sgl_pipe_in(control_sgl_pipe),
    .stop_mark_in(n8091_o),
    .gpr_write_valid_in(gpr_write_valid),
    .gpr_write_in(gpr_write),
    .gpr_a_read_valid_in(gpr_a_read_valid),
    .gpr_a_read_in(gpr_a_read),
    .gpr_b_read_valid_in(gpr_b_read_valid),
    .gpr_b_read_in(gpr_b_read),
    .gpr_c_read_valid_in(gpr_c_read_valid),
    .gpr_c_read_in(gpr_c_read),
    .execute_next_tag_tag(n8093_o),
    .execute_next_tag_valid(n8094_o),
    .execute_next_cr_tag_tag(n8096_o),
    .execute_next_cr_tag_valid(n8097_o),
    .cr_read_in(cr_read_valid),
    .cr_write_in(cr_write_valid),
    .valid_out(control_0_valid_out),
    .stall_out(control_0_stall_out),
    .stopped_out(control_0_stopped_out),
    .gpr_bypass_a(control_0_gpr_bypass_a),
    .gpr_bypass_b(control_0_gpr_bypass_b),
    .gpr_bypass_c(control_0_gpr_bypass_c),
    .cr_bypass(control_0_cr_bypass),
    .instr_tag_out_tag(control_0_instr_tag_out_tag),
    .instr_tag_out_valid(control_0_instr_tag_out_valid));
  assign n8088_o = n8029_o[1:0];
  /* decode1.vhdl:587:44  */
  assign n8089_o = n8029_o[2];
  /* decode2.vhdl:311:30  */
  assign n8090_o = r[392];
  /* decode2.vhdl:316:34  */
  assign n8091_o = n8032_o[1];
  /* decode2.vhdl:330:52  */
  assign n8092_o = n8085_o[2:0];
  /* icache.vhdl:320:14  */
  assign n8093_o = n8092_o[1:0];
  assign n8094_o = n8092_o[2];
  /* decode2.vhdl:331:55  */
  assign n8095_o = n8086_o[2:0];
  /* decode1.vhdl:560:5  */
  assign n8096_o = n8095_o[1:0];
  /* decode1.vhdl:569:18  */
  assign n8097_o = n8095_o[2];
  /* decode1.vhdl:565:18  */
  assign n8105_o = {control_0_instr_tag_out_valid, control_0_instr_tag_out_tag};
  /* decode2.vhdl:348:19  */
  assign n8107_o = r[391:0];
  /* decode2.vhdl:348:21  */
  assign n8108_o = n8107_o[0];
  /* decode2.vhdl:348:27  */
  assign n8109_o = n8108_o & busy_in;
  /* decode2.vhdl:353:26  */
  assign n8112_o = rst | flush_in;
  /* decode2.vhdl:353:56  */
  assign n8113_o = ~deferred;
  /* decode2.vhdl:353:44  */
  assign n8114_o = n8112_o | n8113_o;
  /* decode2.vhdl:362:24  */
  assign n8120_o = n8032_o[162:119];
  /* decode2.vhdl:362:31  */
  assign n8121_o = n8120_o[22];
  assign n8133_o = r[392];
  /* decode2.vhdl:383:31  */
  assign n8134_o = n8032_o[162:119];
  /* decode2.vhdl:383:38  */
  assign n8135_o = n8134_o[23];
  /* decode2.vhdl:386:32  */
  assign n8138_o = n8032_o[162:119];
  /* decode2.vhdl:386:39  */
  assign n8139_o = n8138_o[28];
  assign n8140_o = n8132_o[391:341];
  /* decode2.vhdl:387:19  */
  assign n8141_o = n8032_o[162:119];
  /* decode2.vhdl:387:26  */
  assign n8142_o = n8141_o[8:3];
  /* decode2.vhdl:390:29  */
  assign n8143_o = n8032_o[97:92];
  /* decode2.vhdl:390:44  */
  assign n8145_o = n8143_o == 6'b011111;
  /* decode2.vhdl:390:72  */
  assign n8147_o = n8032_o[97:66];
  /* insn_helpers.vhdl:126:23  */
  assign n8152_o = n8147_o[10];
  /* decode2.vhdl:390:55  */
  assign n8153_o = n8145_o & n8152_o;
  assign n8156_o = n8132_o[331];
  /* decode2.vhdl:390:17  */
  assign n8157_o = n8153_o ? 1'b1 : n8156_o;
  /* decode2.vhdl:390:17  */
  assign n8158_o = n8153_o ? 1'b1 : n8139_o;
  /* decode2.vhdl:388:13  */
  assign n8160_o = n8142_o == 6'b000010;
  /* decode2.vhdl:388:25  */
  assign n8162_o = n8142_o == 6'b101001;
  /* decode2.vhdl:388:25  */
  assign n8163_o = n8160_o | n8162_o;
  /* decode2.vhdl:388:38  */
  assign n8165_o = n8142_o == 6'b010101;
  /* decode2.vhdl:388:38  */
  assign n8166_o = n8163_o | n8165_o;
  /* decode2.vhdl:388:47  */
  assign n8168_o = n8142_o == 6'b010110;
  /* decode2.vhdl:388:47  */
  assign n8169_o = n8166_o | n8168_o;
  /* decode2.vhdl:395:40  */
  assign n8171_o = n8032_o[97:66];
  /* common.vhdl:708:40  */
  assign n8176_o = n8171_o[15:11];
  /* common.vhdl:708:61  */
  assign n8177_o = n8171_o[20:16];
  /* common.vhdl:708:55  */
  assign n8178_o = {n8176_o, n8177_o};
  /* decode2.vhdl:395:46  */
  assign n8180_o = {22'b0, n8178_o};  //  uext
  /* decode2.vhdl:395:46  */
  assign n8182_o = n8180_o == 32'b00000000000000000000000000000001;
  /* decode2.vhdl:395:17  */
  assign n8184_o = n8182_o ? 1'b1 : n8139_o;
  /* decode2.vhdl:394:13  */
  assign n8186_o = n8142_o == 6'b101000;
  assign n8187_o = {n8186_o, n8169_o};
  assign n8188_o = n8132_o[331];
  /* decode2.vhdl:387:9  */
  always @*
    case (n8187_o)
      2'b10: n8189_o = n8188_o;
      2'b01: n8189_o = n8157_o;
      default: n8189_o = n8188_o;
    endcase
  /* decode2.vhdl:387:9  */
  always @*
    case (n8187_o)
      2'b10: n8190_o = n8184_o;
      2'b01: n8190_o = n8158_o;
      default: n8190_o = n8139_o;
    endcase
  assign n8191_o = n8132_o[338:332];
  /* decode2.vhdl:401:51  */
  assign n8194_o = n8032_o[162:119];
  /* decode2.vhdl:401:58  */
  assign n8195_o = n8194_o[11:9];
  /* decode2.vhdl:401:76  */
  assign n8196_o = n8032_o[97:66];
  /* decode2.vhdl:401:87  */
  assign n8197_o = n8074_o[63:0];
  /* decode2.vhdl:401:104  */
  assign n8198_o = n8032_o[104:98];
  /* decode2.vhdl:402:51  */
  assign n8199_o = n8032_o[65:2];
  /* decode2.vhdl:74:14  */
  assign n8205_o = n8195_o == 3'b001;
  /* decode2.vhdl:74:25  */
  assign n8207_o = n8195_o == 3'b010;
  /* insn_helpers.vhdl:61:23  */
  assign n8213_o = n8196_o[20:16];
  /* decode2.vhdl:74:59  */
  assign n8215_o = n8213_o != 5'b00000;
  /* decode2.vhdl:74:38  */
  assign n8216_o = n8207_o & n8215_o;
  /* decode2.vhdl:74:19  */
  assign n8217_o = n8205_o | n8216_o;
  /* insn_helpers.vhdl:61:23  */
  assign n8224_o = n8196_o[20:16];
  /* common.vhdl:761:21  */
  assign n8230_o = {2'b00, n8224_o};
  assign n8232_o = {n8197_o, n8230_o, 1'b1};
  /* decode2.vhdl:76:17  */
  assign n8234_o = n8195_o == 3'b011;
  /* common.vhdl:775:17  */
  assign n8240_o = n8198_o[5];
  assign n8241_o = {n8197_o, n8198_o, n8240_o};
  /* decode2.vhdl:85:17  */
  assign n8243_o = n8195_o == 3'b100;
  assign n8246_o = {n8199_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:87:29  */
  assign n8248_o = n8195_o == 3'b101;
  /* decode2.vhdl:87:23  */
  assign n8250_o = 1'b1 & n8248_o;
  /* insn_helpers.vhdl:236:23  */
  assign n8257_o = n8196_o[20:16];
  /* common.vhdl:780:21  */
  assign n8263_o = {2'b10, n8257_o};
  assign n8265_o = {n8197_o, n8263_o, 1'b1};
  /* decode2.vhdl:87:9  */
  assign n8267_o = n8250_o ? n8265_o : 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
  /* decode2.vhdl:85:9  */
  assign n8268_o = n8243_o ? n8246_o : n8267_o;
  /* decode2.vhdl:76:9  */
  assign n8269_o = n8234_o ? n8241_o : n8268_o;
  /* decode2.vhdl:74:9  */
  assign n8270_o = n8217_o ? n8232_o : n8269_o;
  /* decode2.vhdl:403:51  */
  assign n8272_o = n8032_o[162:119];
  /* decode2.vhdl:403:58  */
  assign n8273_o = n8272_o[15:12];
  /* decode2.vhdl:403:76  */
  assign n8274_o = n8032_o[97:66];
  /* decode2.vhdl:403:87  */
  assign n8275_o = n8074_o[127:64];
  /* decode2.vhdl:403:104  */
  assign n8276_o = n8032_o[111:105];
  /* insn_helpers.vhdl:66:23  */
  assign n8288_o = n8274_o[15:11];
  /* common.vhdl:761:21  */
  assign n8294_o = {2'b00, n8288_o};
  assign n8296_o = {n8275_o, n8294_o, 1'b1};
  /* decode2.vhdl:100:13  */
  assign n8298_o = n8273_o == 4'b0001;
  /* insn_helpers.vhdl:241:23  */
  assign n8305_o = n8274_o[15:11];
  /* common.vhdl:780:21  */
  assign n8311_o = {2'b10, n8305_o};
  assign n8313_o = {n8275_o, n8311_o, 1'b1};
  /* decode2.vhdl:102:13  */
  assign n8315_o = n8273_o == 4'b1111;
  /* insn_helpers.vhdl:81:23  */
  assign n8321_o = n8274_o[15:0];
  /* decode2.vhdl:109:65  */
  assign n8322_o = {48'b0, n8321_o};  //  uext
  assign n8325_o = {n8322_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:108:13  */
  assign n8327_o = n8273_o == 4'b0010;
  /* insn_helpers.vhdl:76:23  */
  assign n8333_o = n8274_o[15:0];
  /* decode2.vhdl:111:65  */
  assign n8334_o = {{48{n8333_o[15]}}, n8333_o}; // sext
  assign n8337_o = {n8334_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:110:13  */
  assign n8339_o = n8273_o == 4'b0011;
  /* insn_helpers.vhdl:76:23  */
  assign n8345_o = n8274_o[15:0];
  /* decode2.vhdl:113:97  */
  assign n8347_o = {n8345_o, 16'b0000000000000000};
  /* decode2.vhdl:113:65  */
  assign n8348_o = {{32{n8347_o[31]}}, n8347_o}; // sext
  assign n8351_o = {n8348_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:112:13  */
  assign n8353_o = n8273_o == 4'b0100;
  /* insn_helpers.vhdl:76:23  */
  assign n8359_o = n8274_o[15:0];
  /* decode2.vhdl:115:99  */
  assign n8361_o = {n8359_o, 16'b0000000000000000};
  /* decode2.vhdl:115:65  */
  assign n8362_o = {32'b0, n8361_o};  //  uext
  assign n8365_o = {n8362_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:114:13  */
  assign n8367_o = n8273_o == 4'b0101;
  /* insn_helpers.vhdl:106:23  */
  assign n8373_o = n8274_o[25:2];
  /* decode2.vhdl:117:97  */
  assign n8375_o = {n8373_o, 2'b00};
  /* decode2.vhdl:117:65  */
  assign n8376_o = {{38{n8375_o[25]}}, n8375_o}; // sext
  assign n8379_o = {n8376_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:116:13  */
  assign n8381_o = n8273_o == 4'b0110;
  /* insn_helpers.vhdl:131:23  */
  assign n8387_o = n8274_o[15:2];
  /* decode2.vhdl:119:97  */
  assign n8389_o = {n8387_o, 2'b00};
  /* decode2.vhdl:119:65  */
  assign n8390_o = {{48{n8389_o[15]}}, n8389_o}; // sext
  assign n8393_o = {n8390_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:118:13  */
  assign n8395_o = n8273_o == 4'b0111;
  /* insn_helpers.vhdl:191:23  */
  assign n8401_o = n8274_o[15:2];
  /* decode2.vhdl:121:97  */
  assign n8403_o = {n8401_o, 2'b00};
  /* decode2.vhdl:121:65  */
  assign n8404_o = {{48{n8403_o[15]}}, n8403_o}; // sext
  assign n8407_o = {n8404_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:120:13  */
  assign n8409_o = n8273_o == 4'b1001;
  /* insn_helpers.vhdl:196:23  */
  assign n8415_o = n8274_o[15:4];
  /* decode2.vhdl:123:97  */
  assign n8417_o = {n8415_o, 4'b0000};
  /* decode2.vhdl:123:65  */
  assign n8418_o = {{48{n8417_o[15]}}, n8417_o}; // sext
  assign n8421_o = {n8418_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:122:13  */
  assign n8423_o = n8273_o == 4'b1010;
  /* insn_helpers.vhdl:201:23  */
  assign n8429_o = n8274_o[15:6];
  /* insn_helpers.vhdl:201:46  */
  assign n8430_o = n8274_o[20:16];
  /* insn_helpers.vhdl:201:37  */
  assign n8431_o = {n8429_o, n8430_o};
  /* insn_helpers.vhdl:201:70  */
  assign n8432_o = n8274_o[0];
  /* insn_helpers.vhdl:201:61  */
  assign n8433_o = {n8431_o, n8432_o};
  /* decode2.vhdl:125:97  */
  assign n8435_o = {n8433_o, 16'b0000000000000100};
  /* decode2.vhdl:125:65  */
  assign n8436_o = {{32{n8435_o[31]}}, n8435_o}; // sext
  assign n8439_o = {n8436_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:124:13  */
  assign n8441_o = n8273_o == 4'b1000;
  /* decode2.vhdl:126:13  */
  assign n8443_o = n8273_o == 4'b1011;
  /* decode2.vhdl:129:81  */
  assign n8444_o = n8274_o[1];
  /* decode2.vhdl:129:72  */
  assign n8446_o = {58'b0000000000000000000000000000000000000000000000000000000000, n8444_o};
  /* decode2.vhdl:129:94  */
  assign n8447_o = n8274_o[15:11];
  /* decode2.vhdl:129:85  */
  assign n8448_o = {n8446_o, n8447_o};
  assign n8451_o = {n8448_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:128:13  */
  assign n8453_o = n8273_o == 4'b1100;
  /* decode2.vhdl:131:82  */
  assign n8454_o = n8274_o[15:11];
  /* decode2.vhdl:131:73  */
  assign n8456_o = {59'b00000000000000000000000000000000000000000000000000000000000, n8454_o};
  assign n8459_o = {n8456_o, 7'b0000000, 1'b0};
  /* decode2.vhdl:130:13  */
  assign n8461_o = n8273_o == 4'b1101;
  /* common.vhdl:775:17  */
  assign n8467_o = n8276_o[5];
  assign n8468_o = {n8275_o, n8276_o, n8467_o};
  /* decode2.vhdl:132:13  */
  assign n8470_o = n8273_o == 4'b1110;
  /* decode2.vhdl:140:13  */
  assign n8472_o = n8273_o == 4'b0000;
  assign n8473_o = {n8472_o, n8470_o, n8461_o, n8453_o, n8443_o, n8441_o, n8423_o, n8409_o, n8395_o, n8381_o, n8367_o, n8353_o, n8339_o, n8327_o, n8315_o, n8298_o};
  /* decode2.vhdl:99:9  */
  always @*
    case (n8473_o)
      16'b1000000000000000: n8477_o = 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
      16'b0100000000000000: n8477_o = n8468_o;
      16'b0010000000000000: n8477_o = n8459_o;
      16'b0001000000000000: n8477_o = n8451_o;
      16'b0000100000000000: n8477_o = 72'b111111111111111111111111111111111111111111111111111111111111111100000000;
      16'b0000010000000000: n8477_o = n8439_o;
      16'b0000001000000000: n8477_o = n8421_o;
      16'b0000000100000000: n8477_o = n8407_o;
      16'b0000000010000000: n8477_o = n8393_o;
      16'b0000000001000000: n8477_o = n8379_o;
      16'b0000000000100000: n8477_o = n8365_o;
      16'b0000000000010000: n8477_o = n8351_o;
      16'b0000000000001000: n8477_o = n8337_o;
      16'b0000000000000100: n8477_o = n8325_o;
      16'b0000000000000010: n8477_o = n8313_o;
      16'b0000000000000001: n8477_o = n8296_o;
      default: n8477_o = 72'bX;
    endcase
  /* decode2.vhdl:404:51  */
  assign n8480_o = n8032_o[162:119];
  /* decode2.vhdl:404:58  */
  assign n8481_o = n8480_o[18:16];
  /* decode2.vhdl:404:76  */
  assign n8482_o = n8032_o[97:66];
  /* decode2.vhdl:404:87  */
  assign n8483_o = n8074_o[191:128];
  /* insn_helpers.vhdl:51:23  */
  assign n8494_o = n8482_o[25:21];
  /* common.vhdl:761:21  */
  assign n8500_o = {2'b00, n8494_o};
  assign n8502_o = {n8483_o, n8500_o, 1'b1};
  /* decode2.vhdl:151:13  */
  assign n8504_o = n8481_o == 3'b001;
  /* insn_helpers.vhdl:71:23  */
  assign n8511_o = n8482_o[10:6];
  /* common.vhdl:761:21  */
  assign n8517_o = {2'b00, n8511_o};
  assign n8519_o = {n8483_o, n8517_o, 1'b1};
  /* decode2.vhdl:153:13  */
  assign n8521_o = n8481_o == 3'b010;
  /* insn_helpers.vhdl:231:23  */
  assign n8528_o = n8482_o[25:21];
  /* common.vhdl:780:21  */
  assign n8534_o = {2'b10, n8528_o};
  assign n8536_o = {n8483_o, n8534_o, 1'b1};
  /* decode2.vhdl:155:13  */
  assign n8538_o = n8481_o == 3'b100;
  /* insn_helpers.vhdl:246:23  */
  assign n8545_o = n8482_o[10:6];
  /* common.vhdl:780:21  */
  assign n8551_o = {2'b10, n8545_o};
  assign n8553_o = {n8483_o, n8551_o, 1'b1};
  /* decode2.vhdl:161:13  */
  assign n8555_o = n8481_o == 3'b011;
  /* decode2.vhdl:167:13  */
  assign n8558_o = n8481_o == 3'b000;
  assign n8559_o = {n8558_o, n8555_o, n8538_o, n8521_o, n8504_o};
  /* decode2.vhdl:150:9  */
  always @*
    case (n8559_o)
      5'b10000: n8561_o = 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
      5'b01000: n8561_o = n8553_o;
      5'b00100: n8561_o = n8536_o;
      5'b00010: n8561_o = n8519_o;
      5'b00001: n8561_o = n8502_o;
      default: n8561_o = 72'bX;
    endcase
  /* decode2.vhdl:405:50  */
  assign n8563_o = n8032_o[162:119];
  /* decode2.vhdl:405:57  */
  assign n8564_o = n8563_o[21:19];
  /* decode2.vhdl:405:76  */
  assign n8565_o = n8032_o[97:66];
  /* decode2.vhdl:405:87  */
  assign n8566_o = n8032_o[118:112];
  /* insn_helpers.vhdl:56:23  */
  assign n8577_o = n8565_o[25:21];
  /* common.vhdl:761:21  */
  assign n8583_o = {2'b00, n8577_o};
  assign n8585_o = {n8583_o, 1'b1};
  /* decode2.vhdl:176:13  */
  assign n8587_o = n8564_o == 3'b001;
  /* insn_helpers.vhdl:61:23  */
  assign n8594_o = n8565_o[20:16];
  /* common.vhdl:761:21  */
  assign n8600_o = {2'b00, n8594_o};
  assign n8602_o = {n8600_o, 1'b1};
  /* decode2.vhdl:178:13  */
  assign n8604_o = n8564_o == 3'b010;
  /* insn_helpers.vhdl:231:23  */
  assign n8611_o = n8565_o[25:21];
  /* common.vhdl:780:21  */
  assign n8617_o = {2'b10, n8611_o};
  assign n8619_o = {n8617_o, 1'b1};
  /* decode2.vhdl:180:13  */
  assign n8621_o = n8564_o == 3'b100;
  /* common.vhdl:775:17  */
  assign n8627_o = n8566_o[5];
  assign n8628_o = {n8566_o, n8627_o};
  /* decode2.vhdl:186:13  */
  assign n8630_o = n8564_o == 3'b011;
  /* decode2.vhdl:194:13  */
  assign n8633_o = n8564_o == 3'b000;
  assign n8634_o = {n8633_o, n8630_o, n8621_o, n8604_o, n8587_o};
  /* decode2.vhdl:175:9  */
  always @*
    case (n8634_o)
      5'b10000: n8636_o = 8'b00000000;
      5'b01000: n8636_o = n8628_o;
      5'b00100: n8636_o = n8619_o;
      5'b00010: n8636_o = n8602_o;
      5'b00001: n8636_o = n8585_o;
      default: n8636_o = 8'bX;
    endcase
  /* decode2.vhdl:407:17  */
  assign n8637_o = n8032_o[162:119];
  /* decode2.vhdl:407:24  */
  assign n8638_o = n8637_o[40];
  /* decode2.vhdl:408:36  */
  assign n8640_o = n8032_o[97:66];
  /* insn_helpers.vhdl:111:23  */
  assign n8645_o = n8640_o[0];
  /* decode2.vhdl:410:40  */
  assign n8647_o = n8032_o[97:66];
  /* insn_helpers.vhdl:116:23  */
  assign n8652_o = n8647_o[1];
  /* decode2.vhdl:410:58  */
  assign n8653_o = n8032_o[92];
  /* decode2.vhdl:410:46  */
  assign n8654_o = n8652_o | n8653_o;
  assign n8655_o = {n8654_o, n8645_o};
  assign n8656_o = n8132_o[329:328];
  /* decode2.vhdl:407:9  */
  assign n8657_o = n8638_o ? n8655_o : n8656_o;
  assign n8658_o = n8132_o[330];
  assign n8659_o = n8132_o[327:0];
  /* decode2.vhdl:412:20  */
  assign n8660_o = n8032_o[162:119];
  /* decode2.vhdl:412:27  */
  assign n8661_o = n8660_o[8:3];
  /* decode2.vhdl:414:17  */
  assign n8662_o = n8032_o[162:119];
  /* decode2.vhdl:414:24  */
  assign n8663_o = n8662_o[43:42];
  /* decode2.vhdl:414:31  */
  assign n8665_o = n8663_o != 2'b00;
  /* decode2.vhdl:416:29  */
  assign n8667_o = r[392];
  /* decode2.vhdl:417:23  */
  assign n8668_o = n8032_o[162:119];
  /* decode2.vhdl:417:30  */
  assign n8669_o = n8668_o[43:42];
  /* decode2.vhdl:420:26  */
  assign n8670_o = r[392];
  /* decode2.vhdl:420:40  */
  assign n8671_o = n8032_o[164];
  /* decode2.vhdl:420:33  */
  assign n8672_o = n8670_o == n8671_o;
  assign n8674_o = n8561_o[1];
  /* decode2.vhdl:420:21  */
  assign n8675_o = n8672_o ? 1'b1 : n8674_o;
  /* decode2.vhdl:418:17  */
  assign n8677_o = n8669_o == 2'b01;
  /* decode2.vhdl:425:26  */
  assign n8678_o = r[392];
  /* decode2.vhdl:425:40  */
  assign n8679_o = n8032_o[164];
  /* decode2.vhdl:425:33  */
  assign n8680_o = n8678_o == n8679_o;
  assign n8682_o = n8636_o[1];
  /* decode2.vhdl:425:21  */
  assign n8683_o = n8680_o ? 1'b1 : n8682_o;
  /* decode2.vhdl:423:17  */
  assign n8685_o = n8669_o == 2'b10;
  /* decode2.vhdl:430:26  */
  assign n8686_o = r[392];
  /* decode2.vhdl:431:60  */
  assign n8687_o = n8270_o[7:1];
  assign n8688_o = n8636_o[7:1];
  /* decode2.vhdl:430:21  */
  assign n8689_o = n8686_o ? n8687_o : n8688_o;
  /* decode2.vhdl:428:17  */
  assign n8691_o = n8669_o == 2'b11;
  assign n8692_o = {n8691_o, n8685_o, n8677_o};
  assign n8693_o = n8561_o[1];
  /* decode2.vhdl:417:13  */
  always @*
    case (n8692_o)
      3'b100: n8694_o = n8693_o;
      3'b010: n8694_o = n8693_o;
      3'b001: n8694_o = n8675_o;
      default: n8694_o = n8693_o;
    endcase
  assign n8695_o = n8689_o[0];
  assign n8696_o = n8636_o[1];
  /* decode2.vhdl:417:13  */
  always @*
    case (n8692_o)
      3'b100: n8697_o = n8695_o;
      3'b010: n8697_o = n8683_o;
      3'b001: n8697_o = n8696_o;
      default: n8697_o = n8696_o;
    endcase
  assign n8698_o = n8689_o[6:1];
  assign n8699_o = n8636_o[7:2];
  /* decode2.vhdl:417:13  */
  always @*
    case (n8692_o)
      3'b100: n8700_o = n8698_o;
      3'b010: n8700_o = n8699_o;
      3'b001: n8700_o = n8699_o;
      default: n8700_o = n8699_o;
    endcase
  assign n8701_o = {n8133_o, n8140_o, n8190_o, n8135_o, n8191_o, n8189_o, n8658_o, n8657_o, n8659_o};
  /* decode2.vhdl:435:17  */
  assign n8702_o = n8701_o[391:0];
  /* decode2.vhdl:435:19  */
  assign n8703_o = n8702_o[328];
  /* decode2.vhdl:435:46  */
  assign n8704_o = n8270_o[0];
  /* decode2.vhdl:435:28  */
  assign n8705_o = n8703_o & n8704_o;
  /* decode2.vhdl:438:29  */
  assign n8707_o = r[392];
  /* decode2.vhdl:440:43  */
  assign n8708_o = r[392];
  /* decode2.vhdl:440:37  */
  assign n8709_o = ~n8708_o;
  assign n8710_o = {n8707_o, 1'b1};
  assign n8711_o = n8132_o[391:390];
  /* decode2.vhdl:435:9  */
  assign n8712_o = n8705_o ? n8710_o : n8711_o;
  assign n8713_o = n8636_o[1];
  /* decode2.vhdl:435:9  */
  assign n8714_o = n8705_o ? n8709_o : n8713_o;
  assign n8715_o = {n8667_o, 1'b1};
  /* decode2.vhdl:414:9  */
  assign n8716_o = n8665_o ? n8715_o : n8712_o;
  assign n8718_o = n8561_o[1];
  /* decode2.vhdl:414:9  */
  assign n8719_o = n8665_o ? n8694_o : n8718_o;
  assign n8720_o = n8561_o[71:2];
  assign n8721_o = n8561_o[0];
  assign n8722_o = {n8700_o, n8697_o};
  assign n8723_o = n8722_o[0];
  /* decode2.vhdl:414:9  */
  assign n8724_o = n8665_o ? n8723_o : n8714_o;
  assign n8725_o = n8722_o[6:1];
  assign n8726_o = n8636_o[7:2];
  /* decode2.vhdl:414:9  */
  assign n8727_o = n8665_o ? n8725_o : n8726_o;
  assign n8729_o = n8636_o[0];
  /* decode2.vhdl:443:45  */
  assign n8730_o = n8270_o[0];
  /* decode2.vhdl:443:64  */
  assign n8731_o = n8032_o[0];
  /* decode2.vhdl:443:55  */
  assign n8732_o = n8730_o & n8731_o;
  /* decode2.vhdl:444:45  */
  assign n8733_o = n8270_o[7:1];
  /* decode2.vhdl:445:45  */
  assign n8734_o = n8477_o[0];
  /* decode2.vhdl:445:64  */
  assign n8735_o = n8032_o[0];
  /* decode2.vhdl:445:55  */
  assign n8736_o = n8734_o & n8735_o;
  /* decode2.vhdl:446:45  */
  assign n8737_o = n8477_o[7:1];
  assign n8738_o = {n8720_o, n8719_o, n8721_o};
  /* decode2.vhdl:447:45  */
  assign n8739_o = n8738_o[0];
  /* decode2.vhdl:447:64  */
  assign n8740_o = n8032_o[0];
  /* decode2.vhdl:447:55  */
  assign n8741_o = n8739_o & n8740_o;
  assign n8742_o = {n8720_o, n8719_o, n8721_o};
  /* decode2.vhdl:448:45  */
  assign n8743_o = n8742_o[7:1];
  /* decode2.vhdl:450:19  */
  assign n8744_o = n8032_o[162:119];
  /* decode2.vhdl:450:26  */
  assign n8745_o = n8744_o[31:29];
  /* decode2.vhdl:451:13  */
  assign n8747_o = n8745_o == 3'b001;
  /* decode2.vhdl:453:13  */
  assign n8749_o = n8745_o == 3'b010;
  /* decode2.vhdl:455:13  */
  assign n8751_o = n8745_o == 3'b011;
  /* decode2.vhdl:457:13  */
  assign n8753_o = n8745_o == 3'b100;
  /* decode2.vhdl:459:13  */
  assign n8755_o = n8745_o == 3'b000;
  assign n8756_o = {n8755_o, n8753_o, n8751_o, n8749_o, n8747_o};
  /* decode2.vhdl:450:9  */
  always @*
    case (n8756_o)
      5'b10000: n8763_o = 4'b0000;
      5'b01000: n8763_o = 4'b1000;
      5'b00100: n8763_o = 4'b0100;
      5'b00010: n8763_o = 4'b0010;
      5'b00001: n8763_o = 4'b0001;
      default: n8763_o = 4'bX;
    endcase
  /* decode2.vhdl:464:25  */
  assign n8764_o = n8032_o[65:2];
  /* decode2.vhdl:465:26  */
  assign n8767_o = n8032_o[162:119];
  /* decode2.vhdl:465:33  */
  assign n8768_o = n8767_o[1:0];
  assign n8770_o = n8132_o[0];
  /* decode2.vhdl:466:25  */
  assign n8771_o = n8032_o[162:119];
  /* decode2.vhdl:466:32  */
  assign n8772_o = n8771_o[2];
  /* decode2.vhdl:468:40  */
  assign n8775_o = n8270_o[7:1];
  /* decode2.vhdl:469:40  */
  assign n8778_o = n8477_o[7:1];
  assign n8780_o = {n8727_o, n8724_o, n8729_o};
  /* decode2.vhdl:470:40  */
  assign n8781_o = n8780_o[7:1];
  assign n8783_o = {n8727_o, n8724_o, n8729_o};
  /* decode2.vhdl:471:47  */
  assign n8784_o = n8783_o[0];
  /* decode2.vhdl:472:34  */
  assign n8786_o = n8032_o[162:119];
  /* decode2.vhdl:472:41  */
  assign n8787_o = n8786_o[39:38];
  /* decode2.vhdl:472:50  */
  assign n8788_o = n8032_o[97:66];
  /* insn_helpers.vhdl:121:23  */
  assign n8798_o = n8788_o[0];
  /* decode2.vhdl:202:13  */
  assign n8800_o = n8787_o == 2'b10;
  /* decode2.vhdl:204:13  */
  assign n8803_o = n8787_o == 2'b01;
  /* decode2.vhdl:206:13  */
  assign n8806_o = n8787_o == 2'b00;
  assign n8807_o = {n8806_o, n8803_o, n8800_o};
  /* decode2.vhdl:201:9  */
  always @*
    case (n8807_o)
      3'b100: n8809_o = 1'b0;
      3'b010: n8809_o = 1'b1;
      3'b001: n8809_o = n8798_o;
      default: n8809_o = 1'bX;
    endcase
  /* decode2.vhdl:473:26  */
  assign n8810_o = n8082_o[36:32];
  /* decode2.vhdl:474:30  */
  assign n8812_o = n8032_o[162:119];
  /* decode2.vhdl:474:37  */
  assign n8813_o = n8812_o[24];
  /* decode2.vhdl:477:32  */
  assign n8817_o = n8032_o[162:119];
  /* decode2.vhdl:477:39  */
  assign n8818_o = n8817_o[25];
  /* decode2.vhdl:478:33  */
  assign n8820_o = n8032_o[162:119];
  /* decode2.vhdl:478:40  */
  assign n8821_o = n8820_o[27:26];
  /* decode2.vhdl:479:34  */
  assign n8823_o = n8032_o[162:119];
  /* decode2.vhdl:479:41  */
  assign n8824_o = n8823_o[28];
  assign n8825_o = n8132_o[338];
  /* decode2.vhdl:480:30  */
  assign n8826_o = n8032_o[162:119];
  /* decode2.vhdl:480:37  */
  assign n8827_o = n8826_o[36];
  /* decode2.vhdl:481:31  */
  assign n8829_o = n8032_o[162:119];
  /* decode2.vhdl:481:38  */
  assign n8830_o = n8829_o[37];
  /* decode2.vhdl:482:26  */
  assign n8832_o = n8032_o[97:66];
  /* decode2.vhdl:484:34  */
  assign n8835_o = n8032_o[162:119];
  /* decode2.vhdl:484:41  */
  assign n8836_o = n8835_o[32];
  /* decode2.vhdl:485:33  */
  assign n8838_o = n8032_o[162:119];
  /* decode2.vhdl:485:40  */
  assign n8839_o = n8838_o[33];
  /* decode2.vhdl:486:28  */
  assign n8841_o = n8032_o[162:119];
  /* decode2.vhdl:486:35  */
  assign n8842_o = n8841_o[34];
  /* decode2.vhdl:487:29  */
  assign n8844_o = n8032_o[162:119];
  /* decode2.vhdl:487:36  */
  assign n8845_o = n8844_o[35];
  /* decode2.vhdl:488:29  */
  assign n8847_o = n8032_o[163];
  /* decode2.vhdl:489:41  */
  assign n8850_o = 6'b111101 - n8661_o;
  /* decode2.vhdl:490:44  */
  assign n8856_o = 6'b111101 - n8661_o;
  /* decode2.vhdl:491:15  */
  assign n8861_o = n8661_o == 6'b000110;
  /* decode2.vhdl:491:29  */
  assign n8863_o = n8661_o == 6'b000111;
  /* decode2.vhdl:491:23  */
  assign n8864_o = n8861_o | n8863_o;
  /* decode2.vhdl:492:25  */
  assign n8865_o = n8032_o[89];
  /* decode2.vhdl:492:30  */
  assign n8866_o = ~n8865_o;
  /* decode2.vhdl:492:42  */
  assign n8867_o = r[392];
  /* decode2.vhdl:492:49  */
  assign n8868_o = ~n8867_o;
  /* decode2.vhdl:492:36  */
  assign n8869_o = n8866_o & n8868_o;
  /* decode2.vhdl:493:27  */
  assign n8870_o = n8032_o[162:119];
  /* decode2.vhdl:493:34  */
  assign n8871_o = n8870_o[8:3];
  /* decode2.vhdl:493:44  */
  assign n8873_o = n8871_o == 6'b000111;
  /* decode2.vhdl:493:68  */
  assign n8874_o = n8032_o[76];
  /* decode2.vhdl:493:73  */
  assign n8875_o = ~n8874_o;
  /* decode2.vhdl:493:55  */
  assign n8876_o = n8873_o & n8875_o;
  /* decode2.vhdl:493:17  */
  assign n8877_o = ~n8876_o;
  /* decode2.vhdl:492:55  */
  assign n8878_o = n8869_o & n8877_o;
  /* decode2.vhdl:491:9  */
  assign n8881_o = n8883_o ? 1'b1 : 1'b0;
  /* decode2.vhdl:491:9  */
  assign n8882_o = n8884_o ? 3'b000 : n8982_data;
  /* decode2.vhdl:491:9  */
  assign n8883_o = n8864_o & n8878_o;
  /* decode2.vhdl:491:9  */
  assign n8884_o = n8864_o & n8878_o;
  /* decode2.vhdl:503:50  */
  assign n8885_o = n8085_o[66:3];
  /* decode2.vhdl:502:13  */
  assign n8887_o = gpr_a_bypass == 1'b1;
  /* decode2.vhdl:505:49  */
  assign n8888_o = n8270_o[71:8];
  /* decode2.vhdl:501:9  */
  always @*
    case (n8887_o)
      1'b1: n8889_o = n8885_o;
      default: n8889_o = n8888_o;
    endcase
  /* decode2.vhdl:509:50  */
  assign n8891_o = n8085_o[66:3];
  /* decode2.vhdl:508:13  */
  assign n8893_o = gpr_b_bypass == 1'b1;
  /* decode2.vhdl:511:49  */
  assign n8894_o = n8477_o[71:8];
  /* decode2.vhdl:507:9  */
  always @*
    case (n8893_o)
      1'b1: n8895_o = n8891_o;
      default: n8895_o = n8894_o;
    endcase
  /* decode2.vhdl:515:50  */
  assign n8897_o = n8085_o[66:3];
  /* decode2.vhdl:514:13  */
  assign n8899_o = gpr_c_bypass == 1'b1;
  assign n8900_o = {n8720_o, n8719_o, n8721_o};
  /* decode2.vhdl:517:49  */
  assign n8901_o = n8900_o[71:8];
  /* decode2.vhdl:513:9  */
  always @*
    case (n8899_o)
      1'b1: n8902_o = n8897_o;
      default: n8902_o = n8901_o;
    endcase
  /* decode2.vhdl:520:24  */
  assign n8904_o = n8082_o[31:0];
  /* decode2.vhdl:522:41  */
  assign n8905_o = n8086_o[34:3];
  /* decode2.vhdl:521:9  */
  assign n8906_o = cr_bypass ? n8905_o : n8904_o;
  /* decode2.vhdl:526:34  */
  assign n8907_o = n8032_o[0];
  /* decode2.vhdl:527:34  */
  assign n8908_o = n8032_o[162:119];
  /* decode2.vhdl:527:41  */
  assign n8909_o = n8908_o[41];
  assign n8910_o = {n8133_o, n8716_o, n8984_data, n8882_o, n8847_o, n8845_o, n8842_o, n8839_o, n8836_o, n8763_o, n8832_o, n8830_o, n8827_o, n8190_o, n8135_o, n8825_o, n8824_o, n8821_o, n8818_o, n8881_o, n8813_o, n8189_o, n8809_o, n8657_o, n8810_o, n8906_o, n8902_o, n8895_o, n8889_o, n8778_o, n8775_o, n8784_o, n8781_o, instr_tag, n8764_o, n8661_o, n8772_o, n8768_o, n8770_o};
  /* decode2.vhdl:529:30  */
  assign n8911_o = n8910_o[391:0];
  /* decode2.vhdl:529:32  */
  assign n8912_o = n8911_o[84];
  assign n8913_o = {n8727_o, n8724_o, n8729_o};
  /* decode2.vhdl:530:36  */
  assign n8914_o = n8913_o[7:1];
  /* decode2.vhdl:532:43  */
  assign n8915_o = n8270_o[0];
  /* decode2.vhdl:533:37  */
  assign n8916_o = n8270_o[7:1];
  /* decode2.vhdl:535:43  */
  assign n8917_o = n8477_o[0];
  /* decode2.vhdl:536:37  */
  assign n8918_o = n8477_o[7:1];
  assign n8919_o = {n8720_o, n8719_o, n8721_o};
  /* decode2.vhdl:538:43  */
  assign n8920_o = n8919_o[0];
  assign n8921_o = {n8720_o, n8719_o, n8721_o};
  /* decode2.vhdl:539:37  */
  assign n8922_o = n8921_o[7:1];
  /* decode2.vhdl:541:32  */
  assign n8923_o = n8032_o[162:119];
  /* decode2.vhdl:541:39  */
  assign n8924_o = n8923_o[23];
  /* decode2.vhdl:541:67  */
  assign n8926_o = n8032_o[162:119];
  /* decode2.vhdl:541:74  */
  assign n8927_o = n8926_o[39:38];
  /* decode2.vhdl:541:83  */
  assign n8928_o = n8032_o[97:66];
  /* insn_helpers.vhdl:121:23  */
  assign n8938_o = n8928_o[0];
  /* decode2.vhdl:202:13  */
  assign n8940_o = n8927_o == 2'b10;
  /* decode2.vhdl:204:13  */
  assign n8943_o = n8927_o == 2'b01;
  /* decode2.vhdl:206:13  */
  assign n8946_o = n8927_o == 2'b00;
  assign n8947_o = {n8946_o, n8943_o, n8940_o};
  /* decode2.vhdl:201:9  */
  always @*
    case (n8947_o)
      3'b100: n8949_o = 1'b0;
      3'b010: n8949_o = 1'b1;
      3'b001: n8949_o = n8938_o;
      default: n8949_o = 1'bX;
    endcase
  /* decode2.vhdl:541:49  */
  assign n8950_o = n8924_o | n8949_o;
  /* decode2.vhdl:544:49  */
  assign n8951_o = n8032_o[162:119];
  /* decode2.vhdl:544:56  */
  assign n8952_o = n8951_o[22];
  /* decode2.vhdl:544:41  */
  assign n8953_o = cr_write_valid | n8952_o;
  assign n8954_o = {n8133_o, n8716_o, n8984_data, n8882_o, n8847_o, n8845_o, n8842_o, n8839_o, n8836_o, n8763_o, n8832_o, n8830_o, n8827_o, n8190_o, n8135_o, n8825_o, n8824_o, n8821_o, n8818_o, n8881_o, n8813_o, n8189_o, n8809_o, n8657_o, n8810_o, n8906_o, n8902_o, n8895_o, n8889_o, n8778_o, n8775_o, n8784_o, n8781_o, instr_tag, n8764_o, n8661_o, n8772_o, n8768_o, control_valid_out};
  /* decode2.vhdl:548:27  */
  assign n8955_o = n8954_o[391:0];
  /* decode2.vhdl:548:29  */
  assign n8956_o = n8955_o[390];
  /* decode2.vhdl:548:46  */
  assign n8957_o = r[392];
  /* decode2.vhdl:548:40  */
  assign n8958_o = ~n8957_o;
  /* decode2.vhdl:548:36  */
  assign n8959_o = n8956_o & n8958_o;
  /* decode2.vhdl:547:9  */
  assign n8960_o = control_valid_out ? n8959_o : n8133_o;
  assign n8961_o = {n8960_o, n8716_o, n8984_data, n8882_o, n8847_o, n8845_o, n8842_o, n8839_o, n8836_o, n8763_o, n8832_o, n8830_o, n8827_o, n8190_o, n8135_o, n8825_o, n8824_o, n8821_o, n8818_o, n8881_o, n8813_o, n8189_o, n8809_o, n8657_o, n8810_o, n8906_o, n8902_o, n8895_o, n8889_o, n8778_o, n8775_o, n8784_o, n8781_o, instr_tag, n8764_o, n8661_o, n8772_o, n8768_o, control_valid_out};
  /* decode2.vhdl:551:45  */
  assign n8962_o = n8961_o[392];
  /* decode2.vhdl:551:40  */
  assign n8963_o = control_stall_out | n8962_o;
  /* decode2.vhdl:553:22  */
  assign n8964_o = rst | flush_in;
  assign n8967_o = {1'b0, 392'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
  assign n8968_o = {n8960_o, n8716_o, n8984_data, n8882_o, n8847_o, n8845_o, n8842_o, n8839_o, n8836_o, n8763_o, n8832_o, n8830_o, n8827_o, n8190_o, n8135_o, n8825_o, n8824_o, n8821_o, n8818_o, n8881_o, n8813_o, n8189_o, n8809_o, n8657_o, n8810_o, n8906_o, n8902_o, n8895_o, n8889_o, n8778_o, n8775_o, n8784_o, n8781_o, instr_tag, n8764_o, n8661_o, n8772_o, n8768_o, control_valid_out};
  /* decode2.vhdl:553:9  */
  assign n8969_o = n8964_o ? n8967_o : n8968_o;
  /* decode2.vhdl:562:20  */
  assign n8970_o = r[391:0];
  /* decode2.vhdl:352:9  */
  assign n8977_o = n8114_o ? rin : r;
  /* decode2.vhdl:352:9  */
  always @(posedge clk)
    n8978_q <= n8977_o;
  /* decode2.vhdl:352:9  */
  assign n8979_o = {n8743_o, n8741_o, n8737_o, n8736_o, n8733_o, n8732_o};
  reg [2:0] n8981[61:0] ; // memory
  initial begin
    n8981[61] = 3'b000;
    n8981[60] = 3'b000;
    n8981[59] = 3'b000;
    n8981[58] = 3'b001;
    n8981[57] = 3'b000;
    n8981[56] = 3'b110;
    n8981[55] = 3'b110;
    n8981[54] = 3'b110;
    n8981[53] = 3'b001;
    n8981[52] = 3'b000;
    n8981[51] = 3'b001;
    n8981[50] = 3'b000;
    n8981[49] = 3'b000;
    n8981[48] = 3'b100;
    n8981[47] = 3'b000;
    n8981[46] = 3'b111;
    n8981[45] = 3'b000;
    n8981[44] = 3'b000;
    n8981[43] = 3'b000;
    n8981[42] = 3'b000;
    n8981[41] = 3'b000;
    n8981[40] = 3'b011;
    n8981[39] = 3'b011;
    n8981[38] = 3'b001;
    n8981[37] = 3'b010;
    n8981[36] = 3'b000;
    n8981[35] = 3'b000;
    n8981[34] = 3'b000;
    n8981[33] = 3'b000;
    n8981[32] = 3'b111;
    n8981[31] = 3'b000;
    n8981[30] = 3'b000;
    n8981[29] = 3'b000;
    n8981[28] = 3'b000;
    n8981[27] = 3'b111;
    n8981[26] = 3'b111;
    n8981[25] = 3'b101;
    n8981[24] = 3'b011;
    n8981[23] = 3'b000;
    n8981[22] = 3'b000;
    n8981[21] = 3'b001;
    n8981[20] = 3'b011;
    n8981[19] = 3'b011;
    n8981[18] = 3'b011;
    n8981[17] = 3'b001;
    n8981[16] = 3'b100;
    n8981[15] = 3'b001;
    n8981[14] = 3'b000;
    n8981[13] = 3'b010;
    n8981[12] = 3'b010;
    n8981[11] = 3'b010;
    n8981[10] = 3'b000;
    n8981[9] = 3'b111;
    n8981[8] = 3'b010;
    n8981[7] = 3'b010;
    n8981[6] = 3'b000;
    n8981[5] = 3'b000;
    n8981[4] = 3'b000;
    n8981[3] = 3'b001;
    n8981[2] = 3'b001;
    n8981[1] = 3'b111;
    n8981[0] = 3'b000;
    end
  assign n8982_data = n8981[n8850_o];
  /* decode2.vhdl:489:41  */
  /* decode2.vhdl:489:40  */
  reg [2:0] n8983[61:0] ; // memory
  initial begin
    n8983[61] = 3'b000;
    n8983[60] = 3'b000;
    n8983[59] = 3'b000;
    n8983[58] = 3'b000;
    n8983[57] = 3'b000;
    n8983[56] = 3'b000;
    n8983[55] = 3'b000;
    n8983[54] = 3'b000;
    n8983[53] = 3'b000;
    n8983[52] = 3'b000;
    n8983[51] = 3'b000;
    n8983[50] = 3'b010;
    n8983[49] = 3'b001;
    n8983[48] = 3'b000;
    n8983[47] = 3'b011;
    n8983[46] = 3'b011;
    n8983[45] = 3'b000;
    n8983[44] = 3'b000;
    n8983[43] = 3'b000;
    n8983[42] = 3'b000;
    n8983[41] = 3'b000;
    n8983[40] = 3'b011;
    n8983[39] = 3'b011;
    n8983[38] = 3'b000;
    n8983[37] = 3'b000;
    n8983[36] = 3'b000;
    n8983[35] = 3'b000;
    n8983[34] = 3'b000;
    n8983[33] = 3'b000;
    n8983[32] = 3'b010;
    n8983[31] = 3'b000;
    n8983[30] = 3'b000;
    n8983[29] = 3'b000;
    n8983[28] = 3'b100;
    n8983[27] = 3'b101;
    n8983[26] = 3'b100;
    n8983[25] = 3'b000;
    n8983[24] = 3'b011;
    n8983[23] = 3'b101;
    n8983[22] = 3'b000;
    n8983[21] = 3'b000;
    n8983[20] = 3'b000;
    n8983[19] = 3'b001;
    n8983[18] = 3'b010;
    n8983[17] = 3'b000;
    n8983[16] = 3'b000;
    n8983[15] = 3'b000;
    n8983[14] = 3'b000;
    n8983[13] = 3'b000;
    n8983[12] = 3'b000;
    n8983[11] = 3'b000;
    n8983[10] = 3'b000;
    n8983[9] = 3'b110;
    n8983[8] = 3'b000;
    n8983[7] = 3'b000;
    n8983[6] = 3'b000;
    n8983[5] = 3'b000;
    n8983[4] = 3'b000;
    n8983[3] = 3'b000;
    n8983[2] = 3'b000;
    n8983[1] = 3'b001;
    n8983[0] = 3'b000;
    end
  assign n8984_data = n8983[n8856_o];
  /* decode2.vhdl:490:44  */
endmodule

module decode1_0_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clk,
   input  rst,
   input  stall_in,
   input  flush_in,
   input  f_in_valid,
   input  f_in_stop_mark,
   input  f_in_fetch_failed,
   input  [63:0] f_in_nia,
   input  [31:0] f_in_insn,
   input  f_in_big_endian,
   input  f_in_next_predicted,
   input  f_in_next_pred_ntaken,
   output busy_out,
   output flush_out,
   output f_out_redirect,
   output [63:0] f_out_redirect_nia,
   output d_out_valid,
   output d_out_stop_mark,
   output [63:0] d_out_nia,
   output [31:0] d_out_insn,
   output [6:0] d_out_ispr1,
   output [6:0] d_out_ispr2,
   output [6:0] d_out_ispro,
   output [43:0] d_out_decode,
   output d_out_br_pred,
   output d_out_big_endian,
   output [12:0] log_out);
  wire [101:0] n7329_o;
  wire n7331_o;
  wire [63:0] n7332_o;
  wire n7334_o;
  wire n7335_o;
  wire [63:0] n7336_o;
  wire [31:0] n7337_o;
  wire [6:0] n7338_o;
  wire [6:0] n7339_o;
  wire [6:0] n7340_o;
  wire [43:0] n7341_o;
  wire n7342_o;
  wire n7343_o;
  wire [164:0] r;
  wire [164:0] rin;
  wire [164:0] s;
  wire [46:0] ri;
  wire [46:0] ri_in;
  wire [46:0] si;
  wire [86:0] br;
  wire [86:0] br_in;
  wire n7349_o;
  wire n7350_o;
  wire [164:0] n7352_o;
  wire n7353_o;
  wire n7354_o;
  wire [46:0] n7355_o;
  wire n7356_o;
  wire n7357_o;
  wire n7358_o;
  wire n7359_o;
  wire [163:0] n7360_o;
  wire n7361_o;
  wire n7362_o;
  wire n7363_o;
  wire n7364_o;
  wire [164:0] n7365_o;
  wire [46:0] n7366_o;
  wire [164:0] n7367_o;
  wire [164:0] n7368_o;
  wire n7369_o;
  wire n7370_o;
  wire [163:0] n7371_o;
  wire [163:0] n7372_o;
  wire [163:0] n7373_o;
  wire [46:0] n7374_o;
  wire [46:0] n7375_o;
  wire n7376_o;
  wire n7377_o;
  wire [163:0] n7378_o;
  wire [163:0] n7379_o;
  wire [163:0] n7380_o;
  wire [164:0] n7381_o;
  wire n7382_o;
  wire n7383_o;
  wire [163:0] n7384_o;
  wire [163:0] n7385_o;
  wire [163:0] n7386_o;
  wire [46:0] n7387_o;
  wire [46:0] n7388_o;
  wire [164:0] n7389_o;
  wire [164:0] n7391_o;
  wire [164:0] n7392_o;
  wire [164:0] n7394_o;
  wire [46:0] n7396_o;
  wire [46:0] n7398_o;
  wire [86:0] n7402_o;
  wire [86:0] n7403_o;
  wire n7410_o;
  wire n7421_o;
  localparam [164:0] n7422_o = 165'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [63:0] n7424_o;
  wire [31:0] n7427_o;
  wire n7429_o;
  wire n7430_o;
  wire [5:0] n7433_o;
  wire [5:0] n7436_o;
  wire n7440_o;
  wire [30:0] n7442_o;
  wire [5:0] n7443_o;
  wire [4:0] n7444_o;
  wire [10:0] n7445_o;
  wire [10:0] n7448_o;
  wire n7452_o;
  wire [5:0] n7453_o;
  wire [5:0] n7456_o;
  wire n7461_o;
  wire [9:0] n7462_o;
  wire [9:0] n7465_o;
  wire [31:0] n7470_o;
  wire [4:0] n7475_o;
  wire [4:0] n7476_o;
  wire [9:0] n7477_o;
  wire n7487_o;
  wire n7489_o;
  wire n7491_o;
  wire n7493_o;
  wire n7495_o;
  wire n7497_o;
  wire n7499_o;
  wire n7501_o;
  wire n7503_o;
  wire n7505_o;
  wire n7507_o;
  wire n7508_o;
  wire n7510_o;
  wire n7512_o;
  wire n7514_o;
  wire n7516_o;
  wire [13:0] n7518_o;
  reg n7521_o;
  reg [6:0] n7527_o;
  reg [4:0] n7543_o;
  wire [4:0] n7547_o;
  wire [6:0] n7550_o;
  wire [6:0] n7555_o;
  wire n7564_o;
  wire n7566_o;
  wire n7568_o;
  wire n7570_o;
  wire n7572_o;
  wire n7574_o;
  wire n7576_o;
  wire n7578_o;
  wire n7580_o;
  wire n7582_o;
  wire n7584_o;
  wire n7585_o;
  wire n7587_o;
  wire n7589_o;
  wire n7591_o;
  wire n7593_o;
  wire [13:0] n7595_o;
  reg n7598_o;
  reg [6:0] n7604_o;
  reg [4:0] n7620_o;
  wire [4:0] n7624_o;
  wire [6:0] n7627_o;
  wire [6:0] n7632_o;
  wire [9:0] n7633_o;
  wire [9:0] n7636_o;
  wire n7637_o;
  wire [6:0] n7639_o;
  wire [164:0] n7640_o;
  wire [6:0] n7641_o;
  wire n7646_o;
  wire n7647_o;
  wire n7652_o;
  wire n7654_o;
  wire n7655_o;
  wire n7657_o;
  wire n7658_o;
  wire n7660_o;
  wire n7661_o;
  reg [1:0] n7663_o;
  reg n7665_o;
  wire [1:0] n7666_o;
  wire [1:0] n7668_o;
  wire [1:0] n7670_o;
  wire [1:0] n7672_o;
  wire [1:0] n7674_o;
  wire [9:0] n7675_o;
  wire [9:0] n7678_o;
  wire n7679_o;
  wire [4:0] n7680_o;
  wire [4:0] n7681_o;
  wire n7682_o;
  wire [4:0] n7683_o;
  wire [4:0] n7684_o;
  wire n7685_o;
  wire n7686_o;
  wire n7689_o;
  wire n7691_o;
  wire n7693_o;
  wire n7694_o;
  wire n7695_o;
  wire n7700_o;
  wire [6:0] n7703_o;
  wire [6:0] n7704_o;
  wire [6:0] n7705_o;
  wire [6:0] n7706_o;
  wire [6:0] n7707_o;
  wire n7708_o;
  wire [13:0] n7709_o;
  wire [23:0] n7710_o;
  wire n7712_o;
  wire [23:0] n7714_o;
  wire n7715_o;
  wire [6:0] n7718_o;
  wire [6:0] n7719_o;
  wire n7721_o;
  wire [4:0] n7722_o;
  wire [4:0] n7723_o;
  wire [9:0] n7724_o;
  wire [9:0] n7727_o;
  wire n7731_o;
  wire n7732_o;
  wire n7733_o;
  wire [1:0] n7734_o;
  wire n7735_o;
  wire [2:0] n7736_o;
  wire [2:0] n7739_o;
  wire n7743_o;
  wire n7744_o;
  wire n7745_o;
  wire n7746_o;
  wire n7747_o;
  wire n7748_o;
  wire n7749_o;
  wire n7750_o;
  wire n7751_o;
  wire n7756_o;
  wire [6:0] n7759_o;
  wire [6:0] n7760_o;
  wire [6:0] n7761_o;
  wire [6:0] n7762_o;
  wire [6:0] n7763_o;
  wire n7764_o;
  wire n7765_o;
  wire n7768_o;
  wire n7769_o;
  wire [6:0] n7774_o;
  wire [6:0] n7775_o;
  wire [13:0] n7780_o;
  wire [20:0] n7781_o;
  wire [13:0] n7782_o;
  wire [13:0] n7783_o;
  wire [6:0] n7784_o;
  wire [6:0] n7785_o;
  wire [6:0] n7786_o;
  wire n7788_o;
  wire [31:0] n7789_o;
  wire [31:0] n7792_o;
  wire n7793_o;
  wire [44:0] n7796_o;
  wire [44:0] n7798_o;
  wire n7800_o;
  wire [3:0] n7801_o;
  wire [3:0] n7804_o;
  wire n7809_o;
  wire [4:0] n7810_o;
  wire [4:0] n7811_o;
  wire n7812_o;
  wire n7815_o;
  wire n7817_o;
  wire [1:0] n7818_o;
  wire [1:0] n7821_o;
  wire n7826_o;
  wire [4:0] n7827_o;
  wire [4:0] n7830_o;
  wire n7834_o;
  wire n7835_o;
  wire [9:0] n7836_o;
  wire [9:0] n7839_o;
  wire n7840_o;
  wire n7841_o;
  wire n7842_o;
  wire n7845_o;
  wire n7847_o;
  wire [1:0] n7848_o;
  wire [1:0] n7851_o;
  wire n7856_o;
  wire n7857_o;
  wire n7858_o;
  wire [3:0] n7859_o;
  wire [4:0] n7860_o;
  wire [8:0] n7861_o;
  wire [8:0] n7864_o;
  wire [3:0] n7868_o;
  wire [4:0] n7870_o;
  wire [4:0] n7872_o;
  wire [43:0] n7876_o;
  wire n7878_o;
  wire [11:0] n7879_o;
  wire [6:0] n7880_o;
  wire [6:0] n7881_o;
  reg [6:0] n7882_o;
  wire [6:0] n7883_o;
  wire [6:0] n7884_o;
  reg [6:0] n7885_o;
  wire [6:0] n7886_o;
  reg [6:0] n7887_o;
  reg [43:0] n7888_o;
  reg n7889_o;
  wire n7892_o;
  reg n7894_o;
  wire [1:0] n7895_o;
  reg [1:0] n7897_o;
  wire [41:0] n7898_o;
  reg [41:0] n7900_o;
  reg [1:0] n7902_o;
  reg [23:0] n7911_o;
  wire n7913_o;
  wire n7917_o;
  wire [43:0] n7918_o;
  wire [5:0] n7919_o;
  wire n7921_o;
  wire n7922_o;
  wire n7924_o;
  wire n7925_o;
  wire [44:0] n7926_o;
  wire [44:0] n7927_o;
  wire [44:0] n7928_o;
  wire [61:0] n7929_o;
  wire n7930_o;
  wire [61:0] n7932_o;
  wire n7933_o;
  wire n7935_o;
  wire n7937_o;
  wire n7938_o;
  wire [164:0] n7939_o;
  wire n7940_o;
  wire n7941_o;
  wire n7942_o;
  wire n7943_o;
  wire n7944_o;
  wire n7945_o;
  wire n7946_o;
  wire n7947_o;
  wire n7948_o;
  wire n7949_o;
  wire [61:0] n7950_o;
  wire [23:0] n7951_o;
  wire [61:0] n7952_o;
  wire [61:0] n7953_o;
  wire [164:0] n7954_o;
  wire [46:0] n7955_o;
  wire [86:0] n7956_o;
  wire n7957_o;
  wire [43:0] n7958_o;
  wire n7959_o;
  wire [43:0] n7960_o;
  wire [1:0] n7961_o;
  wire [1:0] n7962_o;
  wire [1:0] n7963_o;
  wire [1:0] n7964_o;
  wire [1:0] n7965_o;
  wire [118:0] n7970_o;
  wire [1:0] n7971_o;
  wire n7972_o;
  wire n7974_o;
  wire n7975_o;
  wire n7976_o;
  wire n7977_o;
  wire [1:0] n7978_o;
  wire [1:0] n7979_o;
  wire [1:0] n7980_o;
  wire [38:0] n7981_o;
  wire [38:0] n7982_o;
  wire [38:0] n7983_o;
  wire n7984_o;
  wire [63:0] n7986_o;
  wire [86:0] n7987_o;
  wire n7988_o;
  wire n7989_o;
  wire n7990_o;
  reg [164:0] n7995_q;
  reg [164:0] n7996_q;
  reg [46:0] n7999_q;
  reg [46:0] n8000_q;
  reg [86:0] n8001_q;
  wire [64:0] n8002_o;
  wire [164:0] n8003_o;
  localparam [12:0] n8004_o = 13'bZ;
  wire [43:0] n8006_data; // mem_rd
  wire n8008_data; // mem_rd
  wire [43:0] n8010_data; // mem_rd
  wire [43:0] n8012_data; // mem_rd
  wire n8014_data; // mem_rd
  wire [43:0] n8016_data; // mem_rd
  wire [43:0] n8018_data; // mem_rd
  wire [43:0] n8020_data; // mem_rd
  wire [43:0] n8022_data; // mem_rd
  wire [43:0] n8024_data; // mem_rd
  wire [43:0] n8026_data; // mem_rd
  wire [43:0] n8028_data; // mem_rd
  assign busy_out = n7410_o;
  assign flush_out = n7990_o;
  assign f_out_redirect = n7331_o;
  assign f_out_redirect_nia = n7332_o;
  assign d_out_valid = n7334_o;
  assign d_out_stop_mark = n7335_o;
  assign d_out_nia = n7336_o;
  assign d_out_insn = n7337_o;
  assign d_out_ispr1 = n7338_o;
  assign d_out_ispr2 = n7339_o;
  assign d_out_ispro = n7340_o;
  assign d_out_decode = n7341_o;
  assign d_out_br_pred = n7342_o;
  assign d_out_big_endian = n7343_o;
  assign log_out = n8004_o;
  /* icache.vhdl:239:16  */
  assign n7329_o = {f_in_next_pred_ntaken, f_in_next_predicted, f_in_big_endian, f_in_insn, f_in_nia, f_in_fetch_failed, f_in_stop_mark, f_in_valid};
  /* icache.vhdl:237:14  */
  assign n7331_o = n8002_o[0];
  assign n7332_o = n8002_o[64:1];
  assign n7334_o = n8003_o[0];
  assign n7335_o = n8003_o[1];
  /* icache.vhdl:307:14  */
  assign n7336_o = n8003_o[65:2];
  /* icache.vhdl:307:14  */
  assign n7337_o = n8003_o[97:66];
  assign n7338_o = n8003_o[104:98];
  /* icache.vhdl:307:14  */
  assign n7339_o = n8003_o[111:105];
  /* icache.vhdl:301:14  */
  assign n7340_o = n8003_o[118:112];
  /* icache.vhdl:301:14  */
  assign n7341_o = n8003_o[162:119];
  assign n7342_o = n8003_o[163];
  /* icache.vhdl:301:14  */
  assign n7343_o = n8003_o[164];
  /* decode1.vhdl:32:12  */
  assign r = n7995_q; // (signal)
  /* decode1.vhdl:32:15  */
  assign rin = n7954_o; // (signal)
  /* decode1.vhdl:33:12  */
  assign s = n7996_q; // (signal)
  /* decode1.vhdl:48:12  */
  assign ri = n7999_q; // (signal)
  /* decode1.vhdl:48:16  */
  assign ri_in = n7955_o; // (signal)
  /* decode1.vhdl:49:12  */
  assign si = n8000_q; // (signal)
  /* decode1.vhdl:57:12  */
  assign br = n8001_q; // (signal)
  /* decode1.vhdl:57:16  */
  assign br_in = n7956_o; // (signal)
  /* decode1.vhdl:534:21  */
  assign n7349_o = s[0];
  /* decode1.vhdl:535:29  */
  assign n7350_o = ~stall_in;
  /* decode1.vhdl:535:17  */
  assign n7352_o = n7350_o ? s : r;
  /* wishbone_types.vhdl:19:14  */
  assign n7353_o = s[0];
  /* decode1.vhdl:535:17  */
  assign n7354_o = n7350_o ? 1'b0 : n7353_o;
  /* decode1.vhdl:535:17  */
  assign n7355_o = n7350_o ? si : ri;
  /* decode1.vhdl:543:32  */
  assign n7356_o = rin[0];
  /* decode1.vhdl:543:44  */
  assign n7357_o = r[0];
  /* decode1.vhdl:543:38  */
  assign n7358_o = n7356_o & n7357_o;
  /* decode1.vhdl:543:50  */
  assign n7359_o = n7358_o & stall_in;
  /* icache.vhdl:614:18  */
  assign n7360_o = rin[164:1];
  /* decode1.vhdl:544:22  */
  assign n7361_o = r[0];
  /* decode1.vhdl:544:28  */
  assign n7362_o = ~n7361_o;
  /* decode1.vhdl:544:46  */
  assign n7363_o = ~stall_in;
  /* decode1.vhdl:544:34  */
  assign n7364_o = n7362_o | n7363_o;
  /* decode1.vhdl:544:17  */
  assign n7365_o = n7364_o ? rin : r;
  /* decode1.vhdl:544:17  */
  assign n7366_o = n7364_o ? ri_in : ri;
  /* decode1.vhdl:534:13  */
  assign n7367_o = n7349_o ? n7352_o : n7365_o;
  /* icache.vhdl:575:5  */
  assign n7368_o = {n7360_o, n7359_o};
  assign n7369_o = n7368_o[0];
  /* decode1.vhdl:534:13  */
  assign n7370_o = n7349_o ? n7354_o : n7369_o;
  assign n7371_o = n7368_o[164:1];
  /* icache.vhdl:297:43  */
  assign n7372_o = s[164:1];
  /* decode1.vhdl:534:13  */
  assign n7373_o = n7349_o ? n7372_o : n7371_o;
  /* decode1.vhdl:534:13  */
  assign n7374_o = n7349_o ? n7355_o : n7366_o;
  /* decode1.vhdl:534:13  */
  assign n7375_o = n7349_o ? si : ri_in;
  assign n7376_o = n7367_o[0];
  /* decode1.vhdl:531:13  */
  assign n7377_o = flush_in ? 1'b0 : n7376_o;
  assign n7378_o = n7367_o[164:1];
  /* icache.vhdl:297:28  */
  assign n7379_o = r[164:1];
  /* decode1.vhdl:531:13  */
  assign n7380_o = flush_in ? n7379_o : n7378_o;
  /* icache.vhdl:296:17  */
  assign n7381_o = {n7373_o, n7370_o};
  /* icache.vhdl:294:18  */
  assign n7382_o = n7381_o[0];
  /* decode1.vhdl:531:13  */
  assign n7383_o = flush_in ? 1'b0 : n7382_o;
  /* icache.vhdl:292:14  */
  assign n7384_o = n7381_o[164:1];
  /* icache.vhdl:292:14  */
  assign n7385_o = s[164:1];
  /* decode1.vhdl:531:13  */
  assign n7386_o = flush_in ? n7385_o : n7384_o;
  /* decode1.vhdl:531:13  */
  assign n7387_o = flush_in ? ri : n7374_o;
  /* decode1.vhdl:531:13  */
  assign n7388_o = flush_in ? si : n7375_o;
  /* icache.vhdl:545:28  */
  assign n7389_o = {n7380_o, n7377_o};
  /* decode1.vhdl:526:13  */
  assign n7391_o = rst ? 165'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : n7389_o;
  /* icache.vhdl:545:62  */
  assign n7392_o = {n7386_o, n7383_o};
  /* decode1.vhdl:526:13  */
  assign n7394_o = rst ? 165'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : n7392_o;
  /* decode1.vhdl:526:13  */
  assign n7396_o = rst ? 47'b00000000000000000000000000000000000000000000000 : n7387_o;
  /* decode1.vhdl:526:13  */
  assign n7398_o = rst ? 47'b00000000000000000000000000000000000000000000000 : n7388_o;
  /* icache.vhdl:525:40  */
  assign n7402_o = {1'b0, 24'b000000000000000000000000, 62'b00000000000000000000000000000000000000000000000000000000000000};
  /* decode1.vhdl:549:13  */
  assign n7403_o = rst ? n7402_o : br_in;
  /* decode1.vhdl:558:19  */
  assign n7410_o = s[0];
  /* decode1.vhdl:574:25  */
  assign n7421_o = n7329_o[0];
  /* decode1.vhdl:575:24  */
  assign n7424_o = n7329_o[66:3];
  /* decode1.vhdl:576:24  */
  assign n7427_o = n7329_o[98:67];
  /* decode1.vhdl:577:29  */
  assign n7429_o = n7329_o[1];
  /* decode1.vhdl:578:30  */
  assign n7430_o = n7329_o[99];
  /* decode1.vhdl:586:38  */
  assign n7433_o = n7329_o[98:93];
  /* decode1.vhdl:587:44  */
  assign n7436_o = 6'b111111 - n7433_o;
  /* icache.vhdl:320:14  */
  assign n7440_o = n7422_o[163];
  /* decode1.vhdl:589:14  */
  assign n7442_o = {25'b0, n7433_o};  //  uext
  /* decode1.vhdl:592:34  */
  assign n7443_o = n7329_o[72:67];
  /* decode1.vhdl:592:58  */
  assign n7444_o = n7329_o[77:73];
  /* decode1.vhdl:592:47  */
  assign n7445_o = {n7443_o, n7444_o};
  /* decode1.vhdl:593:50  */
  assign n7448_o = 11'b11111111111 - n7445_o;
  /* decode1.vhdl:593:28  */
  assign n7452_o = ~n8008_data;
  /* decode1.vhdl:594:72  */
  assign n7453_o = n7329_o[72:67];
  /* decode1.vhdl:594:43  */
  assign n7456_o = 6'b111111 - n7453_o;
  /* decode1.vhdl:590:9  */
  assign n7461_o = n7442_o == 31'b0000000000000000000000000000100;
  /* decode1.vhdl:598:73  */
  assign n7462_o = n7329_o[77:68];
  /* decode1.vhdl:598:44  */
  assign n7465_o = 10'b1111111111 - n7462_o;
  /* decode1.vhdl:601:41  */
  assign n7470_o = n7329_o[98:67];
  /* common.vhdl:708:40  */
  assign n7475_o = n7470_o[15:11];
  /* common.vhdl:708:61  */
  assign n7476_o = n7470_o[20:16];
  /* common.vhdl:708:55  */
  assign n7477_o = {n7475_o, n7476_o};
  /* common.vhdl:718:8  */
  assign n7487_o = n7477_o == 10'b0000001000;
  /* common.vhdl:720:8  */
  assign n7489_o = n7477_o == 10'b0000001001;
  /* common.vhdl:722:8  */
  assign n7491_o = n7477_o == 10'b0000011010;
  /* common.vhdl:724:8  */
  assign n7493_o = n7477_o == 10'b0000011011;
  /* common.vhdl:726:8  */
  assign n7495_o = n7477_o == 10'b0100111010;
  /* common.vhdl:728:8  */
  assign n7497_o = n7477_o == 10'b0100111011;
  /* common.vhdl:730:8  */
  assign n7499_o = n7477_o == 10'b0100010000;
  /* common.vhdl:732:8  */
  assign n7501_o = n7477_o == 10'b0100010001;
  /* common.vhdl:734:8  */
  assign n7503_o = n7477_o == 10'b0100010010;
  /* common.vhdl:736:8  */
  assign n7505_o = n7477_o == 10'b0100010011;
  /* common.vhdl:736:23  */
  assign n7507_o = n7477_o == 10'b0100000011;
  /* common.vhdl:736:23  */
  assign n7508_o = n7505_o | n7507_o;
  /* common.vhdl:738:8  */
  assign n7510_o = n7477_o == 10'b0100110000;
  /* common.vhdl:740:8  */
  assign n7512_o = n7477_o == 10'b0100110001;
  /* common.vhdl:742:8  */
  assign n7514_o = n7477_o == 10'b0000000001;
  /* common.vhdl:744:8  */
  assign n7516_o = n7477_o == 10'b1100101111;
  assign n7518_o = {n7516_o, n7514_o, n7512_o, n7510_o, n7508_o, n7503_o, n7501_o, n7499_o, n7497_o, n7495_o, n7493_o, n7491_o, n7489_o, n7487_o};
  /* common.vhdl:717:8  */
  always @*
    case (n7518_o)
      14'b10000000000000: n7521_o = 1'b1;
      14'b01000000000000: n7521_o = 1'b1;
      14'b00100000000000: n7521_o = 1'b1;
      14'b00010000000000: n7521_o = 1'b1;
      14'b00001000000000: n7521_o = 1'b1;
      14'b00000100000000: n7521_o = 1'b1;
      14'b00000010000000: n7521_o = 1'b1;
      14'b00000001000000: n7521_o = 1'b1;
      14'b00000000100000: n7521_o = 1'b1;
      14'b00000000010000: n7521_o = 1'b1;
      14'b00000000001000: n7521_o = 1'b1;
      14'b00000000000100: n7521_o = 1'b1;
      14'b00000000000010: n7521_o = 1'b1;
      14'b00000000000001: n7521_o = 1'b1;
      default: n7521_o = 1'b0;
    endcase
  /* common.vhdl:717:8  */
  always @*
    case (n7518_o)
      14'b10000000000000: n7527_o = 7'bX;
      14'b01000000000000: n7527_o = 7'bX;
      14'b00100000000000: n7527_o = 7'bX;
      14'b00010000000000: n7527_o = 7'bX;
      14'b00001000000000: n7527_o = 7'bX;
      14'b00000100000000: n7527_o = 7'bX;
      14'b00000010000000: n7527_o = 7'bX;
      14'b00000001000000: n7527_o = 7'bX;
      14'b00000000100000: n7527_o = 7'bX;
      14'b00000000010000: n7527_o = 7'bX;
      14'b00000000001000: n7527_o = 7'bX;
      14'b00000000000100: n7527_o = 7'bX;
      14'b00000000000010: n7527_o = 7'bX;
      14'b00000000000001: n7527_o = 7'bX;
      default: n7527_o = 7'b0000000;
    endcase
  /* common.vhdl:717:8  */
  always @*
    case (n7518_o)
      14'b10000000000000: n7543_o = 5'b01101;
      14'b01000000000000: n7543_o = 5'b01100;
      14'b00100000000000: n7543_o = 5'b01011;
      14'b00010000000000: n7543_o = 5'b01010;
      14'b00001000000000: n7543_o = 5'b01001;
      14'b00000100000000: n7543_o = 5'b01000;
      14'b00000010000000: n7543_o = 5'b00111;
      14'b00000001000000: n7543_o = 5'b00110;
      14'b00000000100000: n7543_o = 5'b00101;
      14'b00000000010000: n7543_o = 5'b00100;
      14'b00000000001000: n7543_o = 5'b00011;
      14'b00000000000100: n7543_o = 5'b00010;
      14'b00000000000010: n7543_o = 5'b00001;
      14'b00000000000001: n7543_o = 5'b00000;
      default: n7543_o = 5'b00000;
    endcase
  /* common.vhdl:750:8  */
  assign n7547_o = n7521_o ? n7543_o : 5'bXXXXX;
  /* common.vhdl:751:20  */
  assign n7550_o = {2'b01, n7547_o};
  /* common.vhdl:751:8  */
  assign n7555_o = n7521_o ? n7550_o : n7527_o;
  /* common.vhdl:718:8  */
  assign n7564_o = n7477_o == 10'b0000001000;
  /* common.vhdl:720:8  */
  assign n7566_o = n7477_o == 10'b0000001001;
  /* common.vhdl:722:8  */
  assign n7568_o = n7477_o == 10'b0000011010;
  /* common.vhdl:724:8  */
  assign n7570_o = n7477_o == 10'b0000011011;
  /* common.vhdl:726:8  */
  assign n7572_o = n7477_o == 10'b0100111010;
  /* common.vhdl:728:8  */
  assign n7574_o = n7477_o == 10'b0100111011;
  /* common.vhdl:730:8  */
  assign n7576_o = n7477_o == 10'b0100010000;
  /* common.vhdl:732:8  */
  assign n7578_o = n7477_o == 10'b0100010001;
  /* common.vhdl:734:8  */
  assign n7580_o = n7477_o == 10'b0100010010;
  /* common.vhdl:736:8  */
  assign n7582_o = n7477_o == 10'b0100010011;
  /* common.vhdl:736:23  */
  assign n7584_o = n7477_o == 10'b0100000011;
  /* common.vhdl:736:23  */
  assign n7585_o = n7582_o | n7584_o;
  /* common.vhdl:738:8  */
  assign n7587_o = n7477_o == 10'b0100110000;
  /* common.vhdl:740:8  */
  assign n7589_o = n7477_o == 10'b0100110001;
  /* common.vhdl:742:8  */
  assign n7591_o = n7477_o == 10'b0000000001;
  /* common.vhdl:744:8  */
  assign n7593_o = n7477_o == 10'b1100101111;
  assign n7595_o = {n7593_o, n7591_o, n7589_o, n7587_o, n7585_o, n7580_o, n7578_o, n7576_o, n7574_o, n7572_o, n7570_o, n7568_o, n7566_o, n7564_o};
  /* common.vhdl:717:8  */
  always @*
    case (n7595_o)
      14'b10000000000000: n7598_o = 1'b1;
      14'b01000000000000: n7598_o = 1'b1;
      14'b00100000000000: n7598_o = 1'b1;
      14'b00010000000000: n7598_o = 1'b1;
      14'b00001000000000: n7598_o = 1'b1;
      14'b00000100000000: n7598_o = 1'b1;
      14'b00000010000000: n7598_o = 1'b1;
      14'b00000001000000: n7598_o = 1'b1;
      14'b00000000100000: n7598_o = 1'b1;
      14'b00000000010000: n7598_o = 1'b1;
      14'b00000000001000: n7598_o = 1'b1;
      14'b00000000000100: n7598_o = 1'b1;
      14'b00000000000010: n7598_o = 1'b1;
      14'b00000000000001: n7598_o = 1'b1;
      default: n7598_o = 1'b0;
    endcase
  /* common.vhdl:717:8  */
  always @*
    case (n7595_o)
      14'b10000000000000: n7604_o = 7'bX;
      14'b01000000000000: n7604_o = 7'bX;
      14'b00100000000000: n7604_o = 7'bX;
      14'b00010000000000: n7604_o = 7'bX;
      14'b00001000000000: n7604_o = 7'bX;
      14'b00000100000000: n7604_o = 7'bX;
      14'b00000010000000: n7604_o = 7'bX;
      14'b00000001000000: n7604_o = 7'bX;
      14'b00000000100000: n7604_o = 7'bX;
      14'b00000000010000: n7604_o = 7'bX;
      14'b00000000001000: n7604_o = 7'bX;
      14'b00000000000100: n7604_o = 7'bX;
      14'b00000000000010: n7604_o = 7'bX;
      14'b00000000000001: n7604_o = 7'bX;
      default: n7604_o = 7'b0000000;
    endcase
  /* common.vhdl:717:8  */
  always @*
    case (n7595_o)
      14'b10000000000000: n7620_o = 5'b01101;
      14'b01000000000000: n7620_o = 5'b01100;
      14'b00100000000000: n7620_o = 5'b01011;
      14'b00010000000000: n7620_o = 5'b01010;
      14'b00001000000000: n7620_o = 5'b01001;
      14'b00000100000000: n7620_o = 5'b01000;
      14'b00000010000000: n7620_o = 5'b00111;
      14'b00000001000000: n7620_o = 5'b00110;
      14'b00000000100000: n7620_o = 5'b00101;
      14'b00000000010000: n7620_o = 5'b00100;
      14'b00000000001000: n7620_o = 5'b00011;
      14'b00000000000100: n7620_o = 5'b00010;
      14'b00000000000010: n7620_o = 5'b00001;
      14'b00000000000001: n7620_o = 5'b00000;
      default: n7620_o = 5'b00000;
    endcase
  /* common.vhdl:750:8  */
  assign n7624_o = n7598_o ? n7620_o : 5'bXXXXX;
  /* common.vhdl:751:20  */
  assign n7627_o = {2'b01, n7624_o};
  /* common.vhdl:751:8  */
  assign n7632_o = n7598_o ? n7627_o : n7604_o;
  /* decode1.vhdl:605:35  */
  assign n7633_o = n7329_o[77:68];
  /* decode1.vhdl:605:16  */
  assign n7636_o = n7633_o & 10'b1101111111;
  /* decode1.vhdl:605:16  */
  assign n7637_o = n7636_o == 10'b0101010011;
  assign n7639_o = n7422_o[111:105];
  assign n7640_o = {n7430_o, n7440_o, n8012_data, n7632_o, n7639_o, n7555_o, n7427_o, n7424_o, n7429_o, n7421_o};
  /* decode1.vhdl:608:34  */
  assign n7641_o = n7640_o[104:98];
  /* common.vhdl:775:17  */
  assign n7646_o = n7641_o[5];
  /* decode1.vhdl:608:41  */
  assign n7647_o = ~n7646_o;
  /* decode1.vhdl:612:25  */
  assign n7652_o = n7477_o == 10'b0000010011;
  /* decode1.vhdl:612:38  */
  assign n7654_o = n7477_o == 10'b0000010010;
  /* decode1.vhdl:612:38  */
  assign n7655_o = n7652_o | n7654_o;
  /* decode1.vhdl:612:50  */
  assign n7657_o = n7477_o == 10'b0000110000;
  /* decode1.vhdl:612:50  */
  assign n7658_o = n7655_o | n7657_o;
  /* decode1.vhdl:612:60  */
  assign n7660_o = n7477_o == 10'b0111010000;
  /* decode1.vhdl:612:60  */
  assign n7661_o = n7658_o | n7660_o;
  /* decode1.vhdl:611:21  */
  always @*
    case (n7661_o)
      1'b1: n7663_o = 2'b10;
      default: n7663_o = 2'b00;
    endcase
  /* decode1.vhdl:611:21  */
  always @*
    case (n7661_o)
      1'b1: n7665_o = 1'b1;
      default: n7665_o = 1'b0;
    endcase
  assign n7666_o = {1'b1, n7665_o};
  /* decode1.vhdl:608:17  */
  assign n7668_o = n7647_o ? n7663_o : 2'b00;
  /* decode1.vhdl:608:17  */
  assign n7670_o = n7647_o ? n7666_o : 2'b00;
  /* decode1.vhdl:605:13  */
  assign n7672_o = n7637_o ? n7668_o : 2'b00;
  /* decode1.vhdl:605:13  */
  assign n7674_o = n7637_o ? n7670_o : 2'b00;
  /* decode1.vhdl:619:35  */
  assign n7675_o = n7329_o[77:68];
  /* decode1.vhdl:619:16  */
  assign n7678_o = n7675_o & 10'b1111111111;
  /* decode1.vhdl:619:16  */
  assign n7679_o = n7678_o == 10'b0100010100;
  /* decode1.vhdl:621:29  */
  assign n7680_o = n7329_o[92:88];
  /* decode1.vhdl:621:55  */
  assign n7681_o = n7329_o[87:83];
  /* decode1.vhdl:621:44  */
  assign n7682_o = n7680_o == n7681_o;
  /* decode1.vhdl:622:30  */
  assign n7683_o = n7329_o[92:88];
  /* decode1.vhdl:622:56  */
  assign n7684_o = n7329_o[82:78];
  /* decode1.vhdl:622:45  */
  assign n7685_o = n7683_o == n7684_o;
  /* decode1.vhdl:621:70  */
  assign n7686_o = n7682_o | n7685_o;
  /* decode1.vhdl:621:17  */
  assign n7689_o = n7686_o ? 1'b1 : 1'b0;
  /* decode1.vhdl:619:13  */
  assign n7691_o = n7679_o ? n7689_o : 1'b0;
  /* decode1.vhdl:596:9  */
  assign n7693_o = n7442_o == 31'b0000000000000000000000000011111;
  /* decode1.vhdl:629:25  */
  assign n7694_o = n7329_o[90];
  /* decode1.vhdl:629:30  */
  assign n7695_o = ~n7694_o;
  /* decode1.vhdl:632:28  */
  assign n7700_o = n7329_o[67];
  assign n7703_o = n7422_o[118:112];
  /* decode1.vhdl:632:13  */
  assign n7704_o = n7700_o ? 7'b0100000 : n7703_o;
  assign n7705_o = n7422_o[104:98];
  /* decode1.vhdl:629:13  */
  assign n7706_o = n7695_o ? 7'b0100001 : n7705_o;
  /* decode1.vhdl:629:13  */
  assign n7707_o = n7695_o ? 7'b0100001 : n7704_o;
  /* decode1.vhdl:636:35  */
  assign n7708_o = n7329_o[82];
  /* decode1.vhdl:637:49  */
  assign n7709_o = n7329_o[82:69];
  /* decode1.vhdl:637:26  */
  assign n7710_o = {{10{n7709_o[13]}}, n7709_o}; // sext
  /* decode1.vhdl:627:9  */
  assign n7712_o = n7442_o == 31'b0000000000000000000000000010000;
  /* decode1.vhdl:642:42  */
  assign n7714_o = n7329_o[92:69];
  /* decode1.vhdl:643:25  */
  assign n7715_o = n7329_o[67];
  assign n7718_o = n7422_o[118:112];
  /* decode1.vhdl:643:13  */
  assign n7719_o = n7715_o ? 7'b0100000 : n7718_o;
  /* decode1.vhdl:639:9  */
  assign n7721_o = n7442_o == 31'b0000000000000000000000000010010;
  /* decode1.vhdl:648:80  */
  assign n7722_o = n7329_o[72:68];
  /* decode1.vhdl:648:104  */
  assign n7723_o = n7329_o[77:73];
  /* decode1.vhdl:648:93  */
  assign n7724_o = {n7722_o, n7723_o};
  /* decode1.vhdl:648:51  */
  assign n7727_o = 10'b1111111111 - n7724_o;
  /* decode1.vhdl:648:28  */
  assign n7731_o = ~n8014_data;
  /* decode1.vhdl:649:36  */
  assign n7732_o = n7329_o[72];
  /* decode1.vhdl:649:51  */
  assign n7733_o = n7329_o[70];
  /* decode1.vhdl:649:40  */
  assign n7734_o = {n7732_o, n7733_o};
  /* decode1.vhdl:649:66  */
  assign n7735_o = n7329_o[69];
  /* decode1.vhdl:649:55  */
  assign n7736_o = {n7734_o, n7735_o};
  /* decode1.vhdl:650:44  */
  assign n7739_o = 3'b111 - n7736_o;
  /* decode1.vhdl:653:25  */
  assign n7743_o = n7329_o[69];
  /* decode1.vhdl:653:29  */
  assign n7744_o = ~n7743_o;
  /* decode1.vhdl:659:29  */
  assign n7745_o = n7329_o[90];
  /* decode1.vhdl:659:34  */
  assign n7746_o = ~n7745_o;
  /* decode1.vhdl:659:54  */
  assign n7747_o = n7329_o[77];
  /* decode1.vhdl:659:59  */
  assign n7748_o = ~n7747_o;
  /* decode1.vhdl:659:77  */
  assign n7749_o = n7329_o[73];
  /* decode1.vhdl:659:65  */
  assign n7750_o = n7748_o | n7749_o;
  /* decode1.vhdl:659:40  */
  assign n7751_o = n7746_o & n7750_o;
  /* decode1.vhdl:662:32  */
  assign n7756_o = n7329_o[67];
  assign n7759_o = n7422_o[118:112];
  /* decode1.vhdl:662:17  */
  assign n7760_o = n7756_o ? 7'b0100000 : n7759_o;
  assign n7761_o = n7422_o[104:98];
  /* decode1.vhdl:659:17  */
  assign n7762_o = n7751_o ? 7'b0100001 : n7761_o;
  /* decode1.vhdl:659:17  */
  assign n7763_o = n7751_o ? 7'b0100001 : n7760_o;
  /* decode1.vhdl:665:29  */
  assign n7764_o = n7329_o[77];
  /* decode1.vhdl:665:34  */
  assign n7765_o = ~n7764_o;
  /* decode1.vhdl:667:32  */
  assign n7768_o = n7329_o[73];
  /* decode1.vhdl:667:36  */
  assign n7769_o = ~n7768_o;
  /* decode1.vhdl:667:17  */
  assign n7774_o = n7769_o ? 7'b0100001 : 7'b0101101;
  /* decode1.vhdl:665:17  */
  assign n7775_o = n7765_o ? 7'b0100000 : n7774_o;
  assign n7780_o = {7'b0100010, 7'b0100011};
  assign n7781_o = {n7763_o, n7775_o, n7762_o};
  assign n7782_o = n7781_o[13:0];
  /* decode1.vhdl:653:13  */
  assign n7783_o = n7744_o ? n7782_o : n7780_o;
  assign n7784_o = n7781_o[20:14];
  assign n7785_o = n7422_o[118:112];
  /* decode1.vhdl:653:13  */
  assign n7786_o = n7744_o ? n7784_o : n7785_o;
  /* decode1.vhdl:647:9  */
  assign n7788_o = n7442_o == 31'b0000000000000000000000000010011;
  /* decode1.vhdl:680:31  */
  assign n7789_o = n7329_o[98:67];
  /* decode1.vhdl:680:16  */
  assign n7792_o = n7789_o & 32'b11111111111111111111111111111111;
  /* decode1.vhdl:680:16  */
  assign n7793_o = n7792_o == 32'b01100000000000000000000000000000;
  assign n7796_o = {44'b00000000000000000000000000000000000000001001, 1'b1};
  /* decode1.vhdl:680:13  */
  assign n7798_o = n7793_o ? n7796_o : 45'b000000000000000000000000000000000000000000000;
  /* decode1.vhdl:678:9  */
  assign n7800_o = n7442_o == 31'b0000000000000000000000000011000;
  /* decode1.vhdl:687:73  */
  assign n7801_o = n7329_o[71:68];
  /* decode1.vhdl:687:44  */
  assign n7804_o = 4'b1111 - n7801_o;
  /* decode1.vhdl:686:9  */
  assign n7809_o = n7442_o == 31'b0000000000000000000000000011110;
  /* decode1.vhdl:691:25  */
  assign n7810_o = n7329_o[92:88];
  /* decode1.vhdl:691:51  */
  assign n7811_o = n7329_o[87:83];
  /* decode1.vhdl:691:40  */
  assign n7812_o = n7810_o == n7811_o;
  /* decode1.vhdl:691:13  */
  assign n7815_o = n7812_o ? 1'b1 : 1'b0;
  /* decode1.vhdl:689:9  */
  assign n7817_o = n7442_o == 31'b0000000000000000000000000111000;
  /* decode1.vhdl:696:73  */
  assign n7818_o = n7329_o[68:67];
  /* decode1.vhdl:696:44  */
  assign n7821_o = 2'b11 - n7818_o;
  /* decode1.vhdl:695:9  */
  assign n7826_o = n7442_o == 31'b0000000000000000000000000111010;
  /* decode1.vhdl:701:77  */
  assign n7827_o = n7329_o[72:68];
  /* decode1.vhdl:701:48  */
  assign n7830_o = 5'b11111 - n7827_o;
  /* decode1.vhdl:702:29  */
  assign n7834_o = n7329_o[72];
  /* decode1.vhdl:702:33  */
  assign n7835_o = ~n7834_o;
  /* decode1.vhdl:702:66  */
  assign n7836_o = n7329_o[77:68];
  /* decode1.vhdl:702:47  */
  assign n7839_o = n7836_o & 10'b1101111111;
  /* decode1.vhdl:702:47  */
  assign n7840_o = n7839_o == 10'b1101001110;
  /* decode1.vhdl:702:43  */
  assign n7841_o = ~n7840_o;
  /* decode1.vhdl:702:39  */
  assign n7842_o = n7835_o & n7841_o;
  /* decode1.vhdl:702:17  */
  assign n7845_o = n7842_o ? 1'b1 : 1'b0;
  /* decode1.vhdl:698:9  */
  assign n7847_o = n7442_o == 31'b0000000000000000000000000111011;
  /* decode1.vhdl:708:73  */
  assign n7848_o = n7329_o[68:67];
  /* decode1.vhdl:708:44  */
  assign n7851_o = 2'b11 - n7848_o;
  /* decode1.vhdl:707:9  */
  assign n7856_o = n7442_o == 31'b0000000000000000000000000111110;
  /* decode1.vhdl:713:29  */
  assign n7857_o = n7329_o[72];
  /* decode1.vhdl:713:33  */
  assign n7858_o = ~n7857_o;
  /* decode1.vhdl:714:82  */
  assign n7859_o = n7329_o[71:68];
  /* decode1.vhdl:714:106  */
  assign n7860_o = n7329_o[77:73];
  /* decode1.vhdl:714:95  */
  assign n7861_o = {n7859_o, n7860_o};
  /* decode1.vhdl:714:53  */
  assign n7864_o = 9'b111111111 - n7861_o;
  /* decode1.vhdl:716:82  */
  assign n7868_o = n7329_o[71:68];
  /* decode1.vhdl:716:53  */
  assign n7870_o = {1'b0, n7868_o};  //  uext
  /* decode1.vhdl:716:53  */
  assign n7872_o = 5'b10000 - n7870_o;
  /* decode1.vhdl:713:17  */
  assign n7876_o = n7858_o ? n8026_data : n8028_data;
  /* decode1.vhdl:710:9  */
  assign n7878_o = n7442_o == 31'b0000000000000000000000000111111;
  assign n7879_o = {n7878_o, n7856_o, n7847_o, n7826_o, n7817_o, n7809_o, n7800_o, n7788_o, n7721_o, n7712_o, n7693_o, n7461_o};
  assign n7880_o = n7783_o[6:0];
  assign n7881_o = n7422_o[104:98];
  /* decode1.vhdl:589:9  */
  always @*
    case (n7879_o)
      12'b100000000000: n7882_o = n7881_o;
      12'b010000000000: n7882_o = n7881_o;
      12'b001000000000: n7882_o = n7881_o;
      12'b000100000000: n7882_o = n7881_o;
      12'b000010000000: n7882_o = n7881_o;
      12'b000001000000: n7882_o = n7881_o;
      12'b000000100000: n7882_o = n7881_o;
      12'b000000010000: n7882_o = n7880_o;
      12'b000000001000: n7882_o = n7881_o;
      12'b000000000100: n7882_o = n7706_o;
      12'b000000000010: n7882_o = n7555_o;
      12'b000000000001: n7882_o = n7881_o;
      default: n7882_o = n7881_o;
    endcase
  assign n7883_o = n7783_o[13:7];
  assign n7884_o = n7422_o[111:105];
  /* decode1.vhdl:589:9  */
  always @*
    case (n7879_o)
      12'b100000000000: n7885_o = n7884_o;
      12'b010000000000: n7885_o = n7884_o;
      12'b001000000000: n7885_o = n7884_o;
      12'b000100000000: n7885_o = n7884_o;
      12'b000010000000: n7885_o = n7884_o;
      12'b000001000000: n7885_o = n7884_o;
      12'b000000100000: n7885_o = n7884_o;
      12'b000000010000: n7885_o = n7883_o;
      12'b000000001000: n7885_o = n7884_o;
      12'b000000000100: n7885_o = n7884_o;
      12'b000000000010: n7885_o = n7884_o;
      12'b000000000001: n7885_o = n7884_o;
      default: n7885_o = n7884_o;
    endcase
  assign n7886_o = n7422_o[118:112];
  /* decode1.vhdl:589:9  */
  always @*
    case (n7879_o)
      12'b100000000000: n7887_o = n7886_o;
      12'b010000000000: n7887_o = n7886_o;
      12'b001000000000: n7887_o = n7886_o;
      12'b000100000000: n7887_o = n7886_o;
      12'b000010000000: n7887_o = n7886_o;
      12'b000001000000: n7887_o = n7886_o;
      12'b000000100000: n7887_o = n7886_o;
      12'b000000010000: n7887_o = n7786_o;
      12'b000000001000: n7887_o = n7719_o;
      12'b000000000100: n7887_o = n7707_o;
      12'b000000000010: n7887_o = n7632_o;
      12'b000000000001: n7887_o = n7886_o;
      default: n7887_o = n7886_o;
    endcase
  /* decode1.vhdl:589:9  */
  always @*
    case (n7879_o)
      12'b100000000000: n7888_o = n7876_o;
      12'b010000000000: n7888_o = n8024_data;
      12'b001000000000: n7888_o = n8022_data;
      12'b000100000000: n7888_o = n8020_data;
      12'b000010000000: n7888_o = n8006_data;
      12'b000001000000: n7888_o = n8018_data;
      12'b000000100000: n7888_o = n8006_data;
      12'b000000010000: n7888_o = n8016_data;
      12'b000000001000: n7888_o = n8006_data;
      12'b000000000100: n7888_o = n8006_data;
      12'b000000000010: n7888_o = n8012_data;
      12'b000000000001: n7888_o = n8010_data;
      default: n7888_o = n8006_data;
    endcase
  /* decode1.vhdl:589:9  */
  always @*
    case (n7879_o)
      12'b100000000000: n7889_o = n7440_o;
      12'b010000000000: n7889_o = n7440_o;
      12'b001000000000: n7889_o = n7440_o;
      12'b000100000000: n7889_o = n7440_o;
      12'b000010000000: n7889_o = n7440_o;
      12'b000001000000: n7889_o = n7440_o;
      12'b000000100000: n7889_o = n7440_o;
      12'b000000010000: n7889_o = n7440_o;
      12'b000000001000: n7889_o = 1'b1;
      12'b000000000100: n7889_o = n7708_o;
      12'b000000000010: n7889_o = n7440_o;
      12'b000000000001: n7889_o = n7440_o;
      default: n7889_o = n7440_o;
    endcase
  assign n7892_o = n7798_o[0];
  /* decode1.vhdl:589:9  */
  always @*
    case (n7879_o)
      12'b100000000000: n7894_o = 1'b0;
      12'b010000000000: n7894_o = 1'b0;
      12'b001000000000: n7894_o = n7845_o;
      12'b000100000000: n7894_o = 1'b0;
      12'b000010000000: n7894_o = n7815_o;
      12'b000001000000: n7894_o = 1'b0;
      12'b000000100000: n7894_o = n7892_o;
      12'b000000010000: n7894_o = n7731_o;
      12'b000000001000: n7894_o = 1'b0;
      12'b000000000100: n7894_o = 1'b0;
      12'b000000000010: n7894_o = n7691_o;
      12'b000000000001: n7894_o = n7452_o;
      default: n7894_o = 1'b0;
    endcase
  assign n7895_o = n7798_o[2:1];
  /* decode1.vhdl:589:9  */
  always @*
    case (n7879_o)
      12'b100000000000: n7897_o = 2'b00;
      12'b010000000000: n7897_o = 2'b00;
      12'b001000000000: n7897_o = 2'b00;
      12'b000100000000: n7897_o = 2'b00;
      12'b000010000000: n7897_o = 2'b00;
      12'b000001000000: n7897_o = 2'b00;
      12'b000000100000: n7897_o = n7895_o;
      12'b000000010000: n7897_o = 2'b00;
      12'b000000001000: n7897_o = 2'b00;
      12'b000000000100: n7897_o = 2'b00;
      12'b000000000010: n7897_o = n7672_o;
      12'b000000000001: n7897_o = 2'b00;
      default: n7897_o = 2'b00;
    endcase
  assign n7898_o = n7798_o[44:3];
  /* decode1.vhdl:589:9  */
  always @*
    case (n7879_o)
      12'b100000000000: n7900_o = 42'b000000000000000000000000000000000000000000;
      12'b010000000000: n7900_o = 42'b000000000000000000000000000000000000000000;
      12'b001000000000: n7900_o = 42'b000000000000000000000000000000000000000000;
      12'b000100000000: n7900_o = 42'b000000000000000000000000000000000000000000;
      12'b000010000000: n7900_o = 42'b000000000000000000000000000000000000000000;
      12'b000001000000: n7900_o = 42'b000000000000000000000000000000000000000000;
      12'b000000100000: n7900_o = n7898_o;
      12'b000000010000: n7900_o = 42'b000000000000000000000000000000000000000000;
      12'b000000001000: n7900_o = 42'b000000000000000000000000000000000000000000;
      12'b000000000100: n7900_o = 42'b000000000000000000000000000000000000000000;
      12'b000000000010: n7900_o = 42'b000000000000000000000000000000000000000000;
      12'b000000000001: n7900_o = 42'b000000000000000000000000000000000000000000;
      default: n7900_o = 42'b000000000000000000000000000000000000000000;
    endcase
  /* decode1.vhdl:589:9  */
  always @*
    case (n7879_o)
      12'b100000000000: n7902_o = 2'b00;
      12'b010000000000: n7902_o = 2'b00;
      12'b001000000000: n7902_o = 2'b00;
      12'b000100000000: n7902_o = 2'b00;
      12'b000010000000: n7902_o = 2'b00;
      12'b000001000000: n7902_o = 2'b00;
      12'b000000100000: n7902_o = 2'b00;
      12'b000000010000: n7902_o = 2'b00;
      12'b000000001000: n7902_o = 2'b00;
      12'b000000000100: n7902_o = 2'b00;
      12'b000000000010: n7902_o = n7674_o;
      12'b000000000001: n7902_o = 2'b00;
      default: n7902_o = 2'b00;
    endcase
  /* decode1.vhdl:589:9  */
  always @*
    case (n7879_o)
      12'b100000000000: n7911_o = 24'b000000000000000000000000;
      12'b010000000000: n7911_o = 24'b000000000000000000000000;
      12'b001000000000: n7911_o = 24'b000000000000000000000000;
      12'b000100000000: n7911_o = 24'b000000000000000000000000;
      12'b000010000000: n7911_o = 24'b000000000000000000000000;
      12'b000001000000: n7911_o = 24'b000000000000000000000000;
      12'b000000100000: n7911_o = 24'b000000000000000000000000;
      12'b000000010000: n7911_o = 24'b000000000000000000000000;
      12'b000000001000: n7911_o = n7714_o;
      12'b000000000100: n7911_o = n7710_o;
      12'b000000000010: n7911_o = 24'b000000000000000000000000;
      12'b000000000001: n7911_o = 24'b000000000000000000000000;
      default: n7911_o = 24'b000000000000000000000000;
    endcase
  /* decode1.vhdl:723:17  */
  assign n7913_o = n7329_o[2];
  /* decode1.vhdl:728:19  */
  assign n7917_o = ri[0];
  /* decode1.vhdl:728:41  */
  assign n7918_o = ri[44:1];
  /* decode1.vhdl:728:57  */
  assign n7919_o = n7918_o[8:3];
  /* decode1.vhdl:728:67  */
  assign n7921_o = n7919_o == 6'b111101;
  /* decode1.vhdl:728:34  */
  assign n7922_o = n7917_o & n7921_o;
  /* decode1.vhdl:728:13  */
  assign n7924_o = n7922_o ? 1'b0 : 1'b1;
  /* decode1.vhdl:723:9  */
  assign n7925_o = n7913_o ? n7924_o : n7421_o;
  assign n7926_o = {44'b00000000000000000000000000000000000111101010, 1'b1};
  assign n7927_o = {n7900_o, n7897_o, n7894_o};
  /* decode1.vhdl:723:9  */
  assign n7928_o = n7913_o ? n7926_o : n7927_o;
  /* decode1.vhdl:736:30  */
  assign n7929_o = n7329_o[66:5];
  /* decode1.vhdl:737:21  */
  assign n7930_o = n7329_o[68];
  /* decode1.vhdl:737:9  */
  assign n7932_o = n7930_o ? 62'b00000000000000000000000000000000000000000000000000000000000000 : n7929_o;
  /* decode1.vhdl:741:17  */
  assign n7933_o = n7329_o[100];
  /* decode1.vhdl:743:20  */
  assign n7935_o = n7329_o[101];
  /* decode1.vhdl:743:9  */
  assign n7937_o = n7935_o ? 1'b0 : n7889_o;
  /* decode1.vhdl:741:9  */
  assign n7938_o = n7933_o ? 1'b1 : n7937_o;
  assign n7939_o = {n7430_o, n7938_o, n7888_o, n7887_o, n7885_o, n7882_o, n7427_o, n7424_o, n7429_o, n7925_o};
  /* decode1.vhdl:746:25  */
  assign n7940_o = n7939_o[163];
  /* decode1.vhdl:746:42  */
  assign n7941_o = n7329_o[0];
  /* decode1.vhdl:746:33  */
  assign n7942_o = n7940_o & n7941_o;
  /* decode1.vhdl:746:52  */
  assign n7943_o = ~flush_in;
  /* decode1.vhdl:746:48  */
  assign n7944_o = n7942_o & n7943_o;
  /* decode1.vhdl:746:69  */
  assign n7945_o = ~n7410_o;
  /* decode1.vhdl:746:65  */
  assign n7946_o = n7944_o & n7945_o;
  /* decode1.vhdl:746:95  */
  assign n7947_o = n7329_o[100];
  /* decode1.vhdl:746:86  */
  assign n7948_o = ~n7947_o;
  /* decode1.vhdl:746:82  */
  assign n7949_o = n7946_o & n7948_o;
  /* decode1.vhdl:748:50  */
  assign n7950_o = br[61:0];
  /* decode1.vhdl:748:63  */
  assign n7951_o = br[85:62];
  /* decode1.vhdl:748:58  */
  assign n7952_o = {{38{n7951_o[23]}}, n7951_o}; // sext
  /* decode1.vhdl:748:58  */
  assign n7953_o = n7950_o + n7952_o;
  assign n7954_o = {n7430_o, n7938_o, n7888_o, n7887_o, n7885_o, n7882_o, n7427_o, n7424_o, n7429_o, n7925_o};
  assign n7955_o = {n7902_o, n7928_o};
  assign n7956_o = {n7949_o, n7911_o, n7932_o};
  /* decode1.vhdl:757:15  */
  assign n7957_o = ri[0];
  /* decode1.vhdl:758:32  */
  assign n7958_o = ri[44:1];
  /* decode1.vhdl:759:18  */
  assign n7959_o = ri[45];
  /* decode1.vhdl:760:37  */
  assign n7960_o = ri[44:1];
  /* decode1.vhdl:760:53  */
  assign n7961_o = n7960_o[1:0];
  assign n7962_o = r[120:119];
  /* decode1.vhdl:759:9  */
  assign n7963_o = n7959_o ? n7961_o : n7962_o;
  assign n7964_o = n7958_o[1:0];
  /* decode1.vhdl:757:9  */
  assign n7965_o = n7957_o ? n7964_o : n7963_o;
  assign n7970_o = r[118:0];
  assign n7971_o = r[164:163];
  /* decode1.vhdl:762:15  */
  assign n7972_o = ri[46];
  assign n7974_o = ri[42];
  assign n7975_o = r[160];
  /* decode1.vhdl:757:9  */
  assign n7976_o = n7957_o ? n7974_o : n7975_o;
  /* decode1.vhdl:762:9  */
  assign n7977_o = n7972_o ? 1'b1 : n7976_o;
  assign n7978_o = ri[44:43];
  assign n7979_o = r[162:161];
  /* decode1.vhdl:757:9  */
  assign n7980_o = n7957_o ? n7978_o : n7979_o;
  assign n7981_o = ri[41:3];
  assign n7982_o = r[159:121];
  /* decode1.vhdl:757:9  */
  assign n7983_o = n7957_o ? n7981_o : n7982_o;
  /* decode1.vhdl:765:30  */
  assign n7984_o = br[86];
  /* decode1.vhdl:766:41  */
  assign n7986_o = {n7953_o, 2'b00};
  assign n7987_o = {n7949_o, n7911_o, n7932_o};
  /* decode1.vhdl:767:25  */
  assign n7988_o = n7987_o[86];
  /* decode1.vhdl:767:39  */
  assign n7989_o = br[86];
  /* decode1.vhdl:767:33  */
  assign n7990_o = n7988_o | n7989_o;
  /* decode1.vhdl:525:9  */
  always @(posedge clk)
    n7995_q <= n7391_o;
  /* decode1.vhdl:525:9  */
  always @(posedge clk)
    n7996_q <= n7394_o;
  /* decode1.vhdl:525:9  */
  always @(posedge clk)
    n7999_q <= n7396_o;
  /* decode1.vhdl:525:9  */
  always @(posedge clk)
    n8000_q <= n7398_o;
  /* decode1.vhdl:525:9  */
  always @(posedge clk)
    n8001_q <= n7403_o;
  /* decode1.vhdl:525:9  */
  assign n8002_o = {n7986_o, n7984_o};
  assign n8003_o = {n7971_o, n7980_o, n7977_o, n7983_o, n7965_o, n7970_o};
  /* decode1.vhdl:27:9  */
  reg [43:0] n8005[63:0] ; // memory
  initial begin
    n8005[63] = 44'b00100000000000000000000000000000000000100001;
    n8005[62] = 44'b00000000000000000000000000000000000000000000;
    n8005[61] = 44'b00000000000000000000000000000011001111001001;
    n8005[60] = 44'b00000001000000000000000000000011001111001001;
    n8005[59] = 44'b00000000000000000000000000000000000000000000;
    n8005[58] = 44'b00000000000000000000000000000000000000000000;
    n8005[57] = 44'b00000000000000000000000000000000000000000000;
    n8005[56] = 44'b00000010000000000000000010000011001101001001;
    n8005[55] = 44'b00000000000000011101000010000011001000010001;
    n8005[54] = 44'b00000000000000000000000000000000000000000000;
    n8005[53] = 44'b00000000000000001101100000000010001001001001;
    n8005[52] = 44'b00000010000000001101100000000011001001001001;
    n8005[51] = 44'b00000000000000010000000010000011001000010001;
    n8005[50] = 44'b00000100000000010000000010000011001000010001;
    n8005[49] = 44'b00000000000000000000000010000011010000010001;
    n8005[48] = 44'b00000000000000000000000010000100010000010001;
    n8005[47] = 44'b00010000000000000000010110000111011000110001;
    n8005[46] = 44'b00000000000000000000000000000000000110011001;
    n8005[45] = 44'b00010000000000000000000110000110000000101001;
    n8005[44] = 44'b00000000000000000000000000000000000000000000;
    n8005[43] = 44'b00001001000000000000000100011101001110000001;
    n8005[42] = 44'b00001001000000000000000100011101000110000001;
    n8005[41] = 44'b00000000000000000000000000000000000000000000;
    n8005[40] = 44'b00001001000000000000000100010001000110000001;
    n8005[39] = 44'b00000000000000000000000100010010000101100001;
    n8005[38] = 44'b00000000000000000000000100010101000101100001;
    n8005[37] = 44'b00000000000000000000000100010010000111010001;
    n8005[36] = 44'b00000000000000000000000100010101000111010001;
    n8005[35] = 44'b00000100000000000000000100010010000000011001;
    n8005[34] = 44'b00000100000000000000000100010101000000011001;
    n8005[33] = 44'b00000000000000000000000000000000000000000000;
    n8005[32] = 44'b00000000000000000000000000000000000000000000;
    n8005[31] = 44'b00000000000001100000000010000011010011111010;
    n8005[30] = 44'b11000000010001100000000010000011010011111010;
    n8005[29] = 44'b00000000000000100000000010000011010011111010;
    n8005[28] = 44'b11000000010000100000000010000011010011111010;
    n8005[27] = 44'b00000000000001100000000000010011010100000010;
    n8005[26] = 44'b00000000010001100000000100010011010100000010;
    n8005[25] = 44'b00000000000000100000000000010011010100000010;
    n8005[24] = 44'b00000000010000100000000100010011010100000010;
    n8005[23] = 44'b00000000000001000000000010000011010011111010;
    n8005[22] = 44'b11000000010001000000000010000011010011111010;
    n8005[21] = 44'b00000000001001000000000010000011010011111010;
    n8005[20] = 44'b11000000011001000000000010000011010011111010;
    n8005[19] = 44'b00000000000001000000000000010011010100000010;
    n8005[18] = 44'b00000000010001000000000100010011010100000010;
    n8005[17] = 44'b00000000000000000000000000000000000000000000;
    n8005[16] = 44'b00000000000000000000000000000000000000000000;
    n8005[15] = 44'b00000001000001100000001000000011010011111110;
    n8005[14] = 44'b11000001010001100000001000000011010011111110;
    n8005[13] = 44'b00000000000010000000001000000011010011111110;
    n8005[12] = 44'b11000000010010000000001000000011010011111110;
    n8005[11] = 44'b00000001000001100000000001000011010100000110;
    n8005[10] = 44'b00000001010001100000000101000011010100000110;
    n8005[9] = 44'b00000000000010000000000001000011010100000110;
    n8005[8] = 44'b00000000010010000000000101000011010100000110;
    n8005[7] = 44'b10000000000010000000000010001010010011111010;
    n8005[6] = 44'b00000000000000000000000000000000000000000000;
    n8005[5] = 44'b00000000000000000000000000000000000000000000;
    n8005[4] = 44'b00000000000000000000000000000000000000000000;
    n8005[3] = 44'b00000000000000000000000000000000000000000000;
    n8005[2] = 44'b00000000000000000000000000000000000000000000;
    n8005[1] = 44'b00000000000000000000000000000000000000000000;
    n8005[0] = 44'b00000000000000000000000000000000000000000000;
    end
  assign n8006_data = n8005[n7436_o];
  /* decode1.vhdl:587:44  */
  /* decode1.vhdl:587:43  */
  reg n8007[2047:0] ; // memory
  initial begin
    n8007[2047] = 1'b0;
    n8007[2046] = 1'b0;
    n8007[2045] = 1'b0;
    n8007[2044] = 1'b0;
    n8007[2043] = 1'b0;
    n8007[2042] = 1'b0;
    n8007[2041] = 1'b0;
    n8007[2040] = 1'b0;
    n8007[2039] = 1'b0;
    n8007[2038] = 1'b0;
    n8007[2037] = 1'b0;
    n8007[2036] = 1'b0;
    n8007[2035] = 1'b0;
    n8007[2034] = 1'b0;
    n8007[2033] = 1'b0;
    n8007[2032] = 1'b0;
    n8007[2031] = 1'b0;
    n8007[2030] = 1'b0;
    n8007[2029] = 1'b0;
    n8007[2028] = 1'b0;
    n8007[2027] = 1'b0;
    n8007[2026] = 1'b0;
    n8007[2025] = 1'b0;
    n8007[2024] = 1'b0;
    n8007[2023] = 1'b0;
    n8007[2022] = 1'b0;
    n8007[2021] = 1'b0;
    n8007[2020] = 1'b0;
    n8007[2019] = 1'b0;
    n8007[2018] = 1'b0;
    n8007[2017] = 1'b0;
    n8007[2016] = 1'b0;
    n8007[2015] = 1'b0;
    n8007[2014] = 1'b0;
    n8007[2013] = 1'b0;
    n8007[2012] = 1'b0;
    n8007[2011] = 1'b0;
    n8007[2010] = 1'b0;
    n8007[2009] = 1'b0;
    n8007[2008] = 1'b0;
    n8007[2007] = 1'b0;
    n8007[2006] = 1'b0;
    n8007[2005] = 1'b0;
    n8007[2004] = 1'b0;
    n8007[2003] = 1'b0;
    n8007[2002] = 1'b0;
    n8007[2001] = 1'b0;
    n8007[2000] = 1'b0;
    n8007[1999] = 1'b0;
    n8007[1998] = 1'b0;
    n8007[1997] = 1'b0;
    n8007[1996] = 1'b0;
    n8007[1995] = 1'b0;
    n8007[1994] = 1'b0;
    n8007[1993] = 1'b0;
    n8007[1992] = 1'b0;
    n8007[1991] = 1'b0;
    n8007[1990] = 1'b0;
    n8007[1989] = 1'b0;
    n8007[1988] = 1'b0;
    n8007[1987] = 1'b0;
    n8007[1986] = 1'b0;
    n8007[1985] = 1'b0;
    n8007[1984] = 1'b0;
    n8007[1983] = 1'b0;
    n8007[1982] = 1'b0;
    n8007[1981] = 1'b0;
    n8007[1980] = 1'b0;
    n8007[1979] = 1'b0;
    n8007[1978] = 1'b0;
    n8007[1977] = 1'b0;
    n8007[1976] = 1'b0;
    n8007[1975] = 1'b0;
    n8007[1974] = 1'b0;
    n8007[1973] = 1'b0;
    n8007[1972] = 1'b0;
    n8007[1971] = 1'b0;
    n8007[1970] = 1'b0;
    n8007[1969] = 1'b0;
    n8007[1968] = 1'b0;
    n8007[1967] = 1'b0;
    n8007[1966] = 1'b0;
    n8007[1965] = 1'b0;
    n8007[1964] = 1'b0;
    n8007[1963] = 1'b0;
    n8007[1962] = 1'b0;
    n8007[1961] = 1'b0;
    n8007[1960] = 1'b0;
    n8007[1959] = 1'b0;
    n8007[1958] = 1'b0;
    n8007[1957] = 1'b0;
    n8007[1956] = 1'b0;
    n8007[1955] = 1'b0;
    n8007[1954] = 1'b0;
    n8007[1953] = 1'b0;
    n8007[1952] = 1'b0;
    n8007[1951] = 1'b0;
    n8007[1950] = 1'b0;
    n8007[1949] = 1'b0;
    n8007[1948] = 1'b0;
    n8007[1947] = 1'b0;
    n8007[1946] = 1'b0;
    n8007[1945] = 1'b0;
    n8007[1944] = 1'b0;
    n8007[1943] = 1'b0;
    n8007[1942] = 1'b0;
    n8007[1941] = 1'b0;
    n8007[1940] = 1'b0;
    n8007[1939] = 1'b0;
    n8007[1938] = 1'b0;
    n8007[1937] = 1'b0;
    n8007[1936] = 1'b0;
    n8007[1935] = 1'b0;
    n8007[1934] = 1'b0;
    n8007[1933] = 1'b0;
    n8007[1932] = 1'b0;
    n8007[1931] = 1'b0;
    n8007[1930] = 1'b0;
    n8007[1929] = 1'b0;
    n8007[1928] = 1'b0;
    n8007[1927] = 1'b0;
    n8007[1926] = 1'b0;
    n8007[1925] = 1'b0;
    n8007[1924] = 1'b0;
    n8007[1923] = 1'b0;
    n8007[1922] = 1'b0;
    n8007[1921] = 1'b0;
    n8007[1920] = 1'b0;
    n8007[1919] = 1'b0;
    n8007[1918] = 1'b0;
    n8007[1917] = 1'b0;
    n8007[1916] = 1'b0;
    n8007[1915] = 1'b0;
    n8007[1914] = 1'b0;
    n8007[1913] = 1'b0;
    n8007[1912] = 1'b0;
    n8007[1911] = 1'b0;
    n8007[1910] = 1'b0;
    n8007[1909] = 1'b0;
    n8007[1908] = 1'b0;
    n8007[1907] = 1'b0;
    n8007[1906] = 1'b0;
    n8007[1905] = 1'b0;
    n8007[1904] = 1'b0;
    n8007[1903] = 1'b0;
    n8007[1902] = 1'b0;
    n8007[1901] = 1'b0;
    n8007[1900] = 1'b0;
    n8007[1899] = 1'b0;
    n8007[1898] = 1'b0;
    n8007[1897] = 1'b0;
    n8007[1896] = 1'b0;
    n8007[1895] = 1'b0;
    n8007[1894] = 1'b0;
    n8007[1893] = 1'b0;
    n8007[1892] = 1'b0;
    n8007[1891] = 1'b0;
    n8007[1890] = 1'b0;
    n8007[1889] = 1'b0;
    n8007[1888] = 1'b0;
    n8007[1887] = 1'b0;
    n8007[1886] = 1'b0;
    n8007[1885] = 1'b0;
    n8007[1884] = 1'b0;
    n8007[1883] = 1'b0;
    n8007[1882] = 1'b0;
    n8007[1881] = 1'b0;
    n8007[1880] = 1'b0;
    n8007[1879] = 1'b0;
    n8007[1878] = 1'b0;
    n8007[1877] = 1'b0;
    n8007[1876] = 1'b0;
    n8007[1875] = 1'b0;
    n8007[1874] = 1'b0;
    n8007[1873] = 1'b0;
    n8007[1872] = 1'b0;
    n8007[1871] = 1'b0;
    n8007[1870] = 1'b0;
    n8007[1869] = 1'b0;
    n8007[1868] = 1'b0;
    n8007[1867] = 1'b0;
    n8007[1866] = 1'b0;
    n8007[1865] = 1'b0;
    n8007[1864] = 1'b0;
    n8007[1863] = 1'b0;
    n8007[1862] = 1'b0;
    n8007[1861] = 1'b0;
    n8007[1860] = 1'b0;
    n8007[1859] = 1'b0;
    n8007[1858] = 1'b0;
    n8007[1857] = 1'b0;
    n8007[1856] = 1'b0;
    n8007[1855] = 1'b0;
    n8007[1854] = 1'b0;
    n8007[1853] = 1'b0;
    n8007[1852] = 1'b0;
    n8007[1851] = 1'b0;
    n8007[1850] = 1'b0;
    n8007[1849] = 1'b0;
    n8007[1848] = 1'b0;
    n8007[1847] = 1'b0;
    n8007[1846] = 1'b0;
    n8007[1845] = 1'b0;
    n8007[1844] = 1'b0;
    n8007[1843] = 1'b0;
    n8007[1842] = 1'b0;
    n8007[1841] = 1'b0;
    n8007[1840] = 1'b0;
    n8007[1839] = 1'b0;
    n8007[1838] = 1'b0;
    n8007[1837] = 1'b0;
    n8007[1836] = 1'b0;
    n8007[1835] = 1'b0;
    n8007[1834] = 1'b0;
    n8007[1833] = 1'b0;
    n8007[1832] = 1'b0;
    n8007[1831] = 1'b0;
    n8007[1830] = 1'b0;
    n8007[1829] = 1'b0;
    n8007[1828] = 1'b0;
    n8007[1827] = 1'b0;
    n8007[1826] = 1'b0;
    n8007[1825] = 1'b0;
    n8007[1824] = 1'b0;
    n8007[1823] = 1'b0;
    n8007[1822] = 1'b0;
    n8007[1821] = 1'b0;
    n8007[1820] = 1'b0;
    n8007[1819] = 1'b0;
    n8007[1818] = 1'b0;
    n8007[1817] = 1'b0;
    n8007[1816] = 1'b0;
    n8007[1815] = 1'b0;
    n8007[1814] = 1'b0;
    n8007[1813] = 1'b0;
    n8007[1812] = 1'b0;
    n8007[1811] = 1'b0;
    n8007[1810] = 1'b0;
    n8007[1809] = 1'b0;
    n8007[1808] = 1'b0;
    n8007[1807] = 1'b0;
    n8007[1806] = 1'b0;
    n8007[1805] = 1'b0;
    n8007[1804] = 1'b0;
    n8007[1803] = 1'b0;
    n8007[1802] = 1'b0;
    n8007[1801] = 1'b0;
    n8007[1800] = 1'b0;
    n8007[1799] = 1'b0;
    n8007[1798] = 1'b0;
    n8007[1797] = 1'b0;
    n8007[1796] = 1'b0;
    n8007[1795] = 1'b0;
    n8007[1794] = 1'b0;
    n8007[1793] = 1'b0;
    n8007[1792] = 1'b0;
    n8007[1791] = 1'b0;
    n8007[1790] = 1'b0;
    n8007[1789] = 1'b0;
    n8007[1788] = 1'b0;
    n8007[1787] = 1'b0;
    n8007[1786] = 1'b0;
    n8007[1785] = 1'b0;
    n8007[1784] = 1'b0;
    n8007[1783] = 1'b0;
    n8007[1782] = 1'b0;
    n8007[1781] = 1'b0;
    n8007[1780] = 1'b0;
    n8007[1779] = 1'b0;
    n8007[1778] = 1'b0;
    n8007[1777] = 1'b0;
    n8007[1776] = 1'b0;
    n8007[1775] = 1'b0;
    n8007[1774] = 1'b0;
    n8007[1773] = 1'b0;
    n8007[1772] = 1'b0;
    n8007[1771] = 1'b0;
    n8007[1770] = 1'b0;
    n8007[1769] = 1'b0;
    n8007[1768] = 1'b0;
    n8007[1767] = 1'b0;
    n8007[1766] = 1'b0;
    n8007[1765] = 1'b0;
    n8007[1764] = 1'b0;
    n8007[1763] = 1'b0;
    n8007[1762] = 1'b0;
    n8007[1761] = 1'b0;
    n8007[1760] = 1'b0;
    n8007[1759] = 1'b0;
    n8007[1758] = 1'b0;
    n8007[1757] = 1'b0;
    n8007[1756] = 1'b0;
    n8007[1755] = 1'b0;
    n8007[1754] = 1'b0;
    n8007[1753] = 1'b0;
    n8007[1752] = 1'b0;
    n8007[1751] = 1'b0;
    n8007[1750] = 1'b0;
    n8007[1749] = 1'b0;
    n8007[1748] = 1'b0;
    n8007[1747] = 1'b0;
    n8007[1746] = 1'b0;
    n8007[1745] = 1'b0;
    n8007[1744] = 1'b0;
    n8007[1743] = 1'b0;
    n8007[1742] = 1'b0;
    n8007[1741] = 1'b0;
    n8007[1740] = 1'b0;
    n8007[1739] = 1'b0;
    n8007[1738] = 1'b0;
    n8007[1737] = 1'b0;
    n8007[1736] = 1'b0;
    n8007[1735] = 1'b0;
    n8007[1734] = 1'b0;
    n8007[1733] = 1'b0;
    n8007[1732] = 1'b0;
    n8007[1731] = 1'b0;
    n8007[1730] = 1'b0;
    n8007[1729] = 1'b0;
    n8007[1728] = 1'b0;
    n8007[1727] = 1'b0;
    n8007[1726] = 1'b0;
    n8007[1725] = 1'b0;
    n8007[1724] = 1'b0;
    n8007[1723] = 1'b0;
    n8007[1722] = 1'b0;
    n8007[1721] = 1'b0;
    n8007[1720] = 1'b0;
    n8007[1719] = 1'b0;
    n8007[1718] = 1'b0;
    n8007[1717] = 1'b0;
    n8007[1716] = 1'b0;
    n8007[1715] = 1'b0;
    n8007[1714] = 1'b0;
    n8007[1713] = 1'b0;
    n8007[1712] = 1'b0;
    n8007[1711] = 1'b0;
    n8007[1710] = 1'b0;
    n8007[1709] = 1'b0;
    n8007[1708] = 1'b0;
    n8007[1707] = 1'b0;
    n8007[1706] = 1'b0;
    n8007[1705] = 1'b0;
    n8007[1704] = 1'b0;
    n8007[1703] = 1'b0;
    n8007[1702] = 1'b0;
    n8007[1701] = 1'b0;
    n8007[1700] = 1'b0;
    n8007[1699] = 1'b0;
    n8007[1698] = 1'b0;
    n8007[1697] = 1'b0;
    n8007[1696] = 1'b0;
    n8007[1695] = 1'b0;
    n8007[1694] = 1'b0;
    n8007[1693] = 1'b0;
    n8007[1692] = 1'b0;
    n8007[1691] = 1'b0;
    n8007[1690] = 1'b0;
    n8007[1689] = 1'b0;
    n8007[1688] = 1'b0;
    n8007[1687] = 1'b0;
    n8007[1686] = 1'b0;
    n8007[1685] = 1'b0;
    n8007[1684] = 1'b0;
    n8007[1683] = 1'b0;
    n8007[1682] = 1'b0;
    n8007[1681] = 1'b0;
    n8007[1680] = 1'b0;
    n8007[1679] = 1'b0;
    n8007[1678] = 1'b0;
    n8007[1677] = 1'b0;
    n8007[1676] = 1'b0;
    n8007[1675] = 1'b0;
    n8007[1674] = 1'b0;
    n8007[1673] = 1'b0;
    n8007[1672] = 1'b0;
    n8007[1671] = 1'b0;
    n8007[1670] = 1'b0;
    n8007[1669] = 1'b0;
    n8007[1668] = 1'b0;
    n8007[1667] = 1'b0;
    n8007[1666] = 1'b0;
    n8007[1665] = 1'b0;
    n8007[1664] = 1'b0;
    n8007[1663] = 1'b0;
    n8007[1662] = 1'b0;
    n8007[1661] = 1'b0;
    n8007[1660] = 1'b0;
    n8007[1659] = 1'b0;
    n8007[1658] = 1'b0;
    n8007[1657] = 1'b0;
    n8007[1656] = 1'b0;
    n8007[1655] = 1'b0;
    n8007[1654] = 1'b0;
    n8007[1653] = 1'b0;
    n8007[1652] = 1'b0;
    n8007[1651] = 1'b0;
    n8007[1650] = 1'b0;
    n8007[1649] = 1'b0;
    n8007[1648] = 1'b0;
    n8007[1647] = 1'b0;
    n8007[1646] = 1'b0;
    n8007[1645] = 1'b0;
    n8007[1644] = 1'b0;
    n8007[1643] = 1'b0;
    n8007[1642] = 1'b0;
    n8007[1641] = 1'b0;
    n8007[1640] = 1'b0;
    n8007[1639] = 1'b0;
    n8007[1638] = 1'b0;
    n8007[1637] = 1'b0;
    n8007[1636] = 1'b0;
    n8007[1635] = 1'b0;
    n8007[1634] = 1'b0;
    n8007[1633] = 1'b0;
    n8007[1632] = 1'b0;
    n8007[1631] = 1'b0;
    n8007[1630] = 1'b0;
    n8007[1629] = 1'b0;
    n8007[1628] = 1'b0;
    n8007[1627] = 1'b0;
    n8007[1626] = 1'b0;
    n8007[1625] = 1'b0;
    n8007[1624] = 1'b0;
    n8007[1623] = 1'b0;
    n8007[1622] = 1'b0;
    n8007[1621] = 1'b0;
    n8007[1620] = 1'b0;
    n8007[1619] = 1'b0;
    n8007[1618] = 1'b0;
    n8007[1617] = 1'b0;
    n8007[1616] = 1'b0;
    n8007[1615] = 1'b0;
    n8007[1614] = 1'b0;
    n8007[1613] = 1'b0;
    n8007[1612] = 1'b0;
    n8007[1611] = 1'b0;
    n8007[1610] = 1'b0;
    n8007[1609] = 1'b0;
    n8007[1608] = 1'b0;
    n8007[1607] = 1'b0;
    n8007[1606] = 1'b0;
    n8007[1605] = 1'b0;
    n8007[1604] = 1'b0;
    n8007[1603] = 1'b0;
    n8007[1602] = 1'b0;
    n8007[1601] = 1'b0;
    n8007[1600] = 1'b0;
    n8007[1599] = 1'b0;
    n8007[1598] = 1'b0;
    n8007[1597] = 1'b0;
    n8007[1596] = 1'b0;
    n8007[1595] = 1'b0;
    n8007[1594] = 1'b0;
    n8007[1593] = 1'b0;
    n8007[1592] = 1'b0;
    n8007[1591] = 1'b0;
    n8007[1590] = 1'b0;
    n8007[1589] = 1'b0;
    n8007[1588] = 1'b0;
    n8007[1587] = 1'b0;
    n8007[1586] = 1'b0;
    n8007[1585] = 1'b0;
    n8007[1584] = 1'b0;
    n8007[1583] = 1'b0;
    n8007[1582] = 1'b0;
    n8007[1581] = 1'b0;
    n8007[1580] = 1'b0;
    n8007[1579] = 1'b0;
    n8007[1578] = 1'b0;
    n8007[1577] = 1'b0;
    n8007[1576] = 1'b0;
    n8007[1575] = 1'b0;
    n8007[1574] = 1'b0;
    n8007[1573] = 1'b0;
    n8007[1572] = 1'b0;
    n8007[1571] = 1'b0;
    n8007[1570] = 1'b0;
    n8007[1569] = 1'b0;
    n8007[1568] = 1'b0;
    n8007[1567] = 1'b0;
    n8007[1566] = 1'b0;
    n8007[1565] = 1'b0;
    n8007[1564] = 1'b0;
    n8007[1563] = 1'b0;
    n8007[1562] = 1'b0;
    n8007[1561] = 1'b0;
    n8007[1560] = 1'b0;
    n8007[1559] = 1'b0;
    n8007[1558] = 1'b0;
    n8007[1557] = 1'b0;
    n8007[1556] = 1'b0;
    n8007[1555] = 1'b0;
    n8007[1554] = 1'b0;
    n8007[1553] = 1'b0;
    n8007[1552] = 1'b0;
    n8007[1551] = 1'b0;
    n8007[1550] = 1'b0;
    n8007[1549] = 1'b0;
    n8007[1548] = 1'b0;
    n8007[1547] = 1'b0;
    n8007[1546] = 1'b0;
    n8007[1545] = 1'b0;
    n8007[1544] = 1'b0;
    n8007[1543] = 1'b0;
    n8007[1542] = 1'b0;
    n8007[1541] = 1'b0;
    n8007[1540] = 1'b0;
    n8007[1539] = 1'b0;
    n8007[1538] = 1'b0;
    n8007[1537] = 1'b0;
    n8007[1536] = 1'b0;
    n8007[1535] = 1'b0;
    n8007[1534] = 1'b0;
    n8007[1533] = 1'b0;
    n8007[1532] = 1'b0;
    n8007[1531] = 1'b0;
    n8007[1530] = 1'b0;
    n8007[1529] = 1'b0;
    n8007[1528] = 1'b0;
    n8007[1527] = 1'b0;
    n8007[1526] = 1'b0;
    n8007[1525] = 1'b0;
    n8007[1524] = 1'b0;
    n8007[1523] = 1'b0;
    n8007[1522] = 1'b0;
    n8007[1521] = 1'b0;
    n8007[1520] = 1'b0;
    n8007[1519] = 1'b0;
    n8007[1518] = 1'b0;
    n8007[1517] = 1'b0;
    n8007[1516] = 1'b0;
    n8007[1515] = 1'b0;
    n8007[1514] = 1'b0;
    n8007[1513] = 1'b0;
    n8007[1512] = 1'b0;
    n8007[1511] = 1'b0;
    n8007[1510] = 1'b0;
    n8007[1509] = 1'b0;
    n8007[1508] = 1'b0;
    n8007[1507] = 1'b0;
    n8007[1506] = 1'b0;
    n8007[1505] = 1'b0;
    n8007[1504] = 1'b0;
    n8007[1503] = 1'b0;
    n8007[1502] = 1'b0;
    n8007[1501] = 1'b0;
    n8007[1500] = 1'b0;
    n8007[1499] = 1'b0;
    n8007[1498] = 1'b0;
    n8007[1497] = 1'b0;
    n8007[1496] = 1'b0;
    n8007[1495] = 1'b0;
    n8007[1494] = 1'b0;
    n8007[1493] = 1'b0;
    n8007[1492] = 1'b0;
    n8007[1491] = 1'b0;
    n8007[1490] = 1'b0;
    n8007[1489] = 1'b0;
    n8007[1488] = 1'b0;
    n8007[1487] = 1'b0;
    n8007[1486] = 1'b0;
    n8007[1485] = 1'b0;
    n8007[1484] = 1'b0;
    n8007[1483] = 1'b0;
    n8007[1482] = 1'b0;
    n8007[1481] = 1'b0;
    n8007[1480] = 1'b0;
    n8007[1479] = 1'b0;
    n8007[1478] = 1'b0;
    n8007[1477] = 1'b0;
    n8007[1476] = 1'b0;
    n8007[1475] = 1'b0;
    n8007[1474] = 1'b0;
    n8007[1473] = 1'b0;
    n8007[1472] = 1'b0;
    n8007[1471] = 1'b0;
    n8007[1470] = 1'b0;
    n8007[1469] = 1'b0;
    n8007[1468] = 1'b0;
    n8007[1467] = 1'b0;
    n8007[1466] = 1'b0;
    n8007[1465] = 1'b0;
    n8007[1464] = 1'b0;
    n8007[1463] = 1'b0;
    n8007[1462] = 1'b0;
    n8007[1461] = 1'b0;
    n8007[1460] = 1'b0;
    n8007[1459] = 1'b0;
    n8007[1458] = 1'b0;
    n8007[1457] = 1'b0;
    n8007[1456] = 1'b0;
    n8007[1455] = 1'b0;
    n8007[1454] = 1'b0;
    n8007[1453] = 1'b0;
    n8007[1452] = 1'b0;
    n8007[1451] = 1'b0;
    n8007[1450] = 1'b0;
    n8007[1449] = 1'b0;
    n8007[1448] = 1'b0;
    n8007[1447] = 1'b0;
    n8007[1446] = 1'b0;
    n8007[1445] = 1'b0;
    n8007[1444] = 1'b0;
    n8007[1443] = 1'b0;
    n8007[1442] = 1'b0;
    n8007[1441] = 1'b0;
    n8007[1440] = 1'b0;
    n8007[1439] = 1'b0;
    n8007[1438] = 1'b0;
    n8007[1437] = 1'b0;
    n8007[1436] = 1'b0;
    n8007[1435] = 1'b0;
    n8007[1434] = 1'b0;
    n8007[1433] = 1'b0;
    n8007[1432] = 1'b0;
    n8007[1431] = 1'b0;
    n8007[1430] = 1'b0;
    n8007[1429] = 1'b0;
    n8007[1428] = 1'b0;
    n8007[1427] = 1'b0;
    n8007[1426] = 1'b0;
    n8007[1425] = 1'b0;
    n8007[1424] = 1'b0;
    n8007[1423] = 1'b0;
    n8007[1422] = 1'b0;
    n8007[1421] = 1'b0;
    n8007[1420] = 1'b0;
    n8007[1419] = 1'b0;
    n8007[1418] = 1'b0;
    n8007[1417] = 1'b0;
    n8007[1416] = 1'b0;
    n8007[1415] = 1'b0;
    n8007[1414] = 1'b0;
    n8007[1413] = 1'b0;
    n8007[1412] = 1'b0;
    n8007[1411] = 1'b0;
    n8007[1410] = 1'b0;
    n8007[1409] = 1'b0;
    n8007[1408] = 1'b0;
    n8007[1407] = 1'b0;
    n8007[1406] = 1'b0;
    n8007[1405] = 1'b0;
    n8007[1404] = 1'b0;
    n8007[1403] = 1'b0;
    n8007[1402] = 1'b0;
    n8007[1401] = 1'b0;
    n8007[1400] = 1'b0;
    n8007[1399] = 1'b0;
    n8007[1398] = 1'b0;
    n8007[1397] = 1'b0;
    n8007[1396] = 1'b0;
    n8007[1395] = 1'b0;
    n8007[1394] = 1'b0;
    n8007[1393] = 1'b0;
    n8007[1392] = 1'b0;
    n8007[1391] = 1'b0;
    n8007[1390] = 1'b0;
    n8007[1389] = 1'b0;
    n8007[1388] = 1'b0;
    n8007[1387] = 1'b0;
    n8007[1386] = 1'b0;
    n8007[1385] = 1'b0;
    n8007[1384] = 1'b0;
    n8007[1383] = 1'b0;
    n8007[1382] = 1'b0;
    n8007[1381] = 1'b0;
    n8007[1380] = 1'b0;
    n8007[1379] = 1'b0;
    n8007[1378] = 1'b0;
    n8007[1377] = 1'b0;
    n8007[1376] = 1'b0;
    n8007[1375] = 1'b0;
    n8007[1374] = 1'b0;
    n8007[1373] = 1'b0;
    n8007[1372] = 1'b0;
    n8007[1371] = 1'b0;
    n8007[1370] = 1'b0;
    n8007[1369] = 1'b0;
    n8007[1368] = 1'b0;
    n8007[1367] = 1'b0;
    n8007[1366] = 1'b0;
    n8007[1365] = 1'b0;
    n8007[1364] = 1'b0;
    n8007[1363] = 1'b0;
    n8007[1362] = 1'b0;
    n8007[1361] = 1'b0;
    n8007[1360] = 1'b0;
    n8007[1359] = 1'b0;
    n8007[1358] = 1'b0;
    n8007[1357] = 1'b0;
    n8007[1356] = 1'b0;
    n8007[1355] = 1'b0;
    n8007[1354] = 1'b0;
    n8007[1353] = 1'b0;
    n8007[1352] = 1'b0;
    n8007[1351] = 1'b0;
    n8007[1350] = 1'b0;
    n8007[1349] = 1'b0;
    n8007[1348] = 1'b0;
    n8007[1347] = 1'b0;
    n8007[1346] = 1'b0;
    n8007[1345] = 1'b0;
    n8007[1344] = 1'b0;
    n8007[1343] = 1'b0;
    n8007[1342] = 1'b0;
    n8007[1341] = 1'b0;
    n8007[1340] = 1'b0;
    n8007[1339] = 1'b0;
    n8007[1338] = 1'b0;
    n8007[1337] = 1'b0;
    n8007[1336] = 1'b0;
    n8007[1335] = 1'b0;
    n8007[1334] = 1'b0;
    n8007[1333] = 1'b0;
    n8007[1332] = 1'b0;
    n8007[1331] = 1'b0;
    n8007[1330] = 1'b0;
    n8007[1329] = 1'b0;
    n8007[1328] = 1'b0;
    n8007[1327] = 1'b0;
    n8007[1326] = 1'b0;
    n8007[1325] = 1'b0;
    n8007[1324] = 1'b0;
    n8007[1323] = 1'b0;
    n8007[1322] = 1'b0;
    n8007[1321] = 1'b0;
    n8007[1320] = 1'b0;
    n8007[1319] = 1'b0;
    n8007[1318] = 1'b0;
    n8007[1317] = 1'b0;
    n8007[1316] = 1'b0;
    n8007[1315] = 1'b0;
    n8007[1314] = 1'b0;
    n8007[1313] = 1'b0;
    n8007[1312] = 1'b0;
    n8007[1311] = 1'b0;
    n8007[1310] = 1'b0;
    n8007[1309] = 1'b0;
    n8007[1308] = 1'b0;
    n8007[1307] = 1'b0;
    n8007[1306] = 1'b0;
    n8007[1305] = 1'b0;
    n8007[1304] = 1'b0;
    n8007[1303] = 1'b0;
    n8007[1302] = 1'b0;
    n8007[1301] = 1'b0;
    n8007[1300] = 1'b0;
    n8007[1299] = 1'b0;
    n8007[1298] = 1'b0;
    n8007[1297] = 1'b0;
    n8007[1296] = 1'b0;
    n8007[1295] = 1'b0;
    n8007[1294] = 1'b0;
    n8007[1293] = 1'b0;
    n8007[1292] = 1'b0;
    n8007[1291] = 1'b0;
    n8007[1290] = 1'b0;
    n8007[1289] = 1'b0;
    n8007[1288] = 1'b0;
    n8007[1287] = 1'b0;
    n8007[1286] = 1'b0;
    n8007[1285] = 1'b0;
    n8007[1284] = 1'b0;
    n8007[1283] = 1'b0;
    n8007[1282] = 1'b0;
    n8007[1281] = 1'b0;
    n8007[1280] = 1'b0;
    n8007[1279] = 1'b0;
    n8007[1278] = 1'b0;
    n8007[1277] = 1'b0;
    n8007[1276] = 1'b0;
    n8007[1275] = 1'b0;
    n8007[1274] = 1'b0;
    n8007[1273] = 1'b0;
    n8007[1272] = 1'b0;
    n8007[1271] = 1'b0;
    n8007[1270] = 1'b0;
    n8007[1269] = 1'b0;
    n8007[1268] = 1'b0;
    n8007[1267] = 1'b0;
    n8007[1266] = 1'b0;
    n8007[1265] = 1'b0;
    n8007[1264] = 1'b0;
    n8007[1263] = 1'b0;
    n8007[1262] = 1'b0;
    n8007[1261] = 1'b0;
    n8007[1260] = 1'b0;
    n8007[1259] = 1'b0;
    n8007[1258] = 1'b0;
    n8007[1257] = 1'b0;
    n8007[1256] = 1'b0;
    n8007[1255] = 1'b0;
    n8007[1254] = 1'b0;
    n8007[1253] = 1'b0;
    n8007[1252] = 1'b0;
    n8007[1251] = 1'b0;
    n8007[1250] = 1'b0;
    n8007[1249] = 1'b0;
    n8007[1248] = 1'b0;
    n8007[1247] = 1'b0;
    n8007[1246] = 1'b0;
    n8007[1245] = 1'b0;
    n8007[1244] = 1'b0;
    n8007[1243] = 1'b0;
    n8007[1242] = 1'b0;
    n8007[1241] = 1'b0;
    n8007[1240] = 1'b0;
    n8007[1239] = 1'b0;
    n8007[1238] = 1'b0;
    n8007[1237] = 1'b0;
    n8007[1236] = 1'b0;
    n8007[1235] = 1'b0;
    n8007[1234] = 1'b0;
    n8007[1233] = 1'b0;
    n8007[1232] = 1'b0;
    n8007[1231] = 1'b0;
    n8007[1230] = 1'b0;
    n8007[1229] = 1'b0;
    n8007[1228] = 1'b0;
    n8007[1227] = 1'b0;
    n8007[1226] = 1'b0;
    n8007[1225] = 1'b0;
    n8007[1224] = 1'b0;
    n8007[1223] = 1'b0;
    n8007[1222] = 1'b0;
    n8007[1221] = 1'b0;
    n8007[1220] = 1'b0;
    n8007[1219] = 1'b0;
    n8007[1218] = 1'b0;
    n8007[1217] = 1'b0;
    n8007[1216] = 1'b0;
    n8007[1215] = 1'b0;
    n8007[1214] = 1'b0;
    n8007[1213] = 1'b0;
    n8007[1212] = 1'b0;
    n8007[1211] = 1'b0;
    n8007[1210] = 1'b0;
    n8007[1209] = 1'b0;
    n8007[1208] = 1'b0;
    n8007[1207] = 1'b0;
    n8007[1206] = 1'b0;
    n8007[1205] = 1'b0;
    n8007[1204] = 1'b0;
    n8007[1203] = 1'b0;
    n8007[1202] = 1'b0;
    n8007[1201] = 1'b0;
    n8007[1200] = 1'b0;
    n8007[1199] = 1'b0;
    n8007[1198] = 1'b0;
    n8007[1197] = 1'b0;
    n8007[1196] = 1'b0;
    n8007[1195] = 1'b0;
    n8007[1194] = 1'b0;
    n8007[1193] = 1'b0;
    n8007[1192] = 1'b0;
    n8007[1191] = 1'b0;
    n8007[1190] = 1'b0;
    n8007[1189] = 1'b0;
    n8007[1188] = 1'b0;
    n8007[1187] = 1'b0;
    n8007[1186] = 1'b0;
    n8007[1185] = 1'b0;
    n8007[1184] = 1'b0;
    n8007[1183] = 1'b0;
    n8007[1182] = 1'b0;
    n8007[1181] = 1'b0;
    n8007[1180] = 1'b0;
    n8007[1179] = 1'b0;
    n8007[1178] = 1'b0;
    n8007[1177] = 1'b0;
    n8007[1176] = 1'b0;
    n8007[1175] = 1'b0;
    n8007[1174] = 1'b0;
    n8007[1173] = 1'b0;
    n8007[1172] = 1'b0;
    n8007[1171] = 1'b0;
    n8007[1170] = 1'b0;
    n8007[1169] = 1'b0;
    n8007[1168] = 1'b0;
    n8007[1167] = 1'b0;
    n8007[1166] = 1'b0;
    n8007[1165] = 1'b0;
    n8007[1164] = 1'b0;
    n8007[1163] = 1'b0;
    n8007[1162] = 1'b0;
    n8007[1161] = 1'b0;
    n8007[1160] = 1'b0;
    n8007[1159] = 1'b0;
    n8007[1158] = 1'b0;
    n8007[1157] = 1'b0;
    n8007[1156] = 1'b0;
    n8007[1155] = 1'b0;
    n8007[1154] = 1'b0;
    n8007[1153] = 1'b0;
    n8007[1152] = 1'b0;
    n8007[1151] = 1'b0;
    n8007[1150] = 1'b0;
    n8007[1149] = 1'b0;
    n8007[1148] = 1'b0;
    n8007[1147] = 1'b0;
    n8007[1146] = 1'b0;
    n8007[1145] = 1'b0;
    n8007[1144] = 1'b0;
    n8007[1143] = 1'b0;
    n8007[1142] = 1'b0;
    n8007[1141] = 1'b0;
    n8007[1140] = 1'b0;
    n8007[1139] = 1'b0;
    n8007[1138] = 1'b0;
    n8007[1137] = 1'b0;
    n8007[1136] = 1'b0;
    n8007[1135] = 1'b0;
    n8007[1134] = 1'b0;
    n8007[1133] = 1'b0;
    n8007[1132] = 1'b0;
    n8007[1131] = 1'b0;
    n8007[1130] = 1'b0;
    n8007[1129] = 1'b0;
    n8007[1128] = 1'b0;
    n8007[1127] = 1'b0;
    n8007[1126] = 1'b0;
    n8007[1125] = 1'b0;
    n8007[1124] = 1'b0;
    n8007[1123] = 1'b0;
    n8007[1122] = 1'b0;
    n8007[1121] = 1'b0;
    n8007[1120] = 1'b0;
    n8007[1119] = 1'b0;
    n8007[1118] = 1'b0;
    n8007[1117] = 1'b0;
    n8007[1116] = 1'b0;
    n8007[1115] = 1'b0;
    n8007[1114] = 1'b0;
    n8007[1113] = 1'b0;
    n8007[1112] = 1'b0;
    n8007[1111] = 1'b0;
    n8007[1110] = 1'b0;
    n8007[1109] = 1'b0;
    n8007[1108] = 1'b0;
    n8007[1107] = 1'b0;
    n8007[1106] = 1'b0;
    n8007[1105] = 1'b0;
    n8007[1104] = 1'b0;
    n8007[1103] = 1'b0;
    n8007[1102] = 1'b0;
    n8007[1101] = 1'b0;
    n8007[1100] = 1'b0;
    n8007[1099] = 1'b0;
    n8007[1098] = 1'b0;
    n8007[1097] = 1'b0;
    n8007[1096] = 1'b0;
    n8007[1095] = 1'b0;
    n8007[1094] = 1'b0;
    n8007[1093] = 1'b0;
    n8007[1092] = 1'b0;
    n8007[1091] = 1'b0;
    n8007[1090] = 1'b0;
    n8007[1089] = 1'b0;
    n8007[1088] = 1'b0;
    n8007[1087] = 1'b0;
    n8007[1086] = 1'b0;
    n8007[1085] = 1'b0;
    n8007[1084] = 1'b0;
    n8007[1083] = 1'b0;
    n8007[1082] = 1'b0;
    n8007[1081] = 1'b0;
    n8007[1080] = 1'b0;
    n8007[1079] = 1'b0;
    n8007[1078] = 1'b0;
    n8007[1077] = 1'b0;
    n8007[1076] = 1'b0;
    n8007[1075] = 1'b0;
    n8007[1074] = 1'b0;
    n8007[1073] = 1'b0;
    n8007[1072] = 1'b0;
    n8007[1071] = 1'b0;
    n8007[1070] = 1'b0;
    n8007[1069] = 1'b0;
    n8007[1068] = 1'b0;
    n8007[1067] = 1'b0;
    n8007[1066] = 1'b0;
    n8007[1065] = 1'b0;
    n8007[1064] = 1'b0;
    n8007[1063] = 1'b0;
    n8007[1062] = 1'b0;
    n8007[1061] = 1'b0;
    n8007[1060] = 1'b0;
    n8007[1059] = 1'b0;
    n8007[1058] = 1'b0;
    n8007[1057] = 1'b0;
    n8007[1056] = 1'b0;
    n8007[1055] = 1'b0;
    n8007[1054] = 1'b0;
    n8007[1053] = 1'b0;
    n8007[1052] = 1'b0;
    n8007[1051] = 1'b0;
    n8007[1050] = 1'b0;
    n8007[1049] = 1'b0;
    n8007[1048] = 1'b0;
    n8007[1047] = 1'b0;
    n8007[1046] = 1'b0;
    n8007[1045] = 1'b0;
    n8007[1044] = 1'b0;
    n8007[1043] = 1'b0;
    n8007[1042] = 1'b0;
    n8007[1041] = 1'b0;
    n8007[1040] = 1'b0;
    n8007[1039] = 1'b0;
    n8007[1038] = 1'b0;
    n8007[1037] = 1'b0;
    n8007[1036] = 1'b0;
    n8007[1035] = 1'b0;
    n8007[1034] = 1'b0;
    n8007[1033] = 1'b0;
    n8007[1032] = 1'b0;
    n8007[1031] = 1'b0;
    n8007[1030] = 1'b0;
    n8007[1029] = 1'b0;
    n8007[1028] = 1'b0;
    n8007[1027] = 1'b0;
    n8007[1026] = 1'b0;
    n8007[1025] = 1'b0;
    n8007[1024] = 1'b0;
    n8007[1023] = 1'b0;
    n8007[1022] = 1'b0;
    n8007[1021] = 1'b0;
    n8007[1020] = 1'b0;
    n8007[1019] = 1'b0;
    n8007[1018] = 1'b0;
    n8007[1017] = 1'b0;
    n8007[1016] = 1'b0;
    n8007[1015] = 1'b0;
    n8007[1014] = 1'b0;
    n8007[1013] = 1'b0;
    n8007[1012] = 1'b0;
    n8007[1011] = 1'b0;
    n8007[1010] = 1'b0;
    n8007[1009] = 1'b0;
    n8007[1008] = 1'b0;
    n8007[1007] = 1'b0;
    n8007[1006] = 1'b0;
    n8007[1005] = 1'b0;
    n8007[1004] = 1'b0;
    n8007[1003] = 1'b0;
    n8007[1002] = 1'b0;
    n8007[1001] = 1'b0;
    n8007[1000] = 1'b0;
    n8007[999] = 1'b0;
    n8007[998] = 1'b0;
    n8007[997] = 1'b0;
    n8007[996] = 1'b0;
    n8007[995] = 1'b0;
    n8007[994] = 1'b0;
    n8007[993] = 1'b0;
    n8007[992] = 1'b0;
    n8007[991] = 1'b0;
    n8007[990] = 1'b0;
    n8007[989] = 1'b0;
    n8007[988] = 1'b0;
    n8007[987] = 1'b0;
    n8007[986] = 1'b0;
    n8007[985] = 1'b0;
    n8007[984] = 1'b0;
    n8007[983] = 1'b0;
    n8007[982] = 1'b0;
    n8007[981] = 1'b0;
    n8007[980] = 1'b0;
    n8007[979] = 1'b0;
    n8007[978] = 1'b0;
    n8007[977] = 1'b0;
    n8007[976] = 1'b0;
    n8007[975] = 1'b0;
    n8007[974] = 1'b0;
    n8007[973] = 1'b0;
    n8007[972] = 1'b0;
    n8007[971] = 1'b0;
    n8007[970] = 1'b0;
    n8007[969] = 1'b0;
    n8007[968] = 1'b0;
    n8007[967] = 1'b0;
    n8007[966] = 1'b0;
    n8007[965] = 1'b0;
    n8007[964] = 1'b0;
    n8007[963] = 1'b0;
    n8007[962] = 1'b0;
    n8007[961] = 1'b0;
    n8007[960] = 1'b0;
    n8007[959] = 1'b0;
    n8007[958] = 1'b0;
    n8007[957] = 1'b0;
    n8007[956] = 1'b0;
    n8007[955] = 1'b0;
    n8007[954] = 1'b0;
    n8007[953] = 1'b0;
    n8007[952] = 1'b0;
    n8007[951] = 1'b0;
    n8007[950] = 1'b0;
    n8007[949] = 1'b0;
    n8007[948] = 1'b0;
    n8007[947] = 1'b0;
    n8007[946] = 1'b0;
    n8007[945] = 1'b0;
    n8007[944] = 1'b0;
    n8007[943] = 1'b0;
    n8007[942] = 1'b0;
    n8007[941] = 1'b0;
    n8007[940] = 1'b0;
    n8007[939] = 1'b0;
    n8007[938] = 1'b0;
    n8007[937] = 1'b0;
    n8007[936] = 1'b0;
    n8007[935] = 1'b0;
    n8007[934] = 1'b0;
    n8007[933] = 1'b0;
    n8007[932] = 1'b0;
    n8007[931] = 1'b0;
    n8007[930] = 1'b0;
    n8007[929] = 1'b0;
    n8007[928] = 1'b0;
    n8007[927] = 1'b0;
    n8007[926] = 1'b0;
    n8007[925] = 1'b0;
    n8007[924] = 1'b0;
    n8007[923] = 1'b0;
    n8007[922] = 1'b0;
    n8007[921] = 1'b0;
    n8007[920] = 1'b0;
    n8007[919] = 1'b0;
    n8007[918] = 1'b0;
    n8007[917] = 1'b0;
    n8007[916] = 1'b0;
    n8007[915] = 1'b0;
    n8007[914] = 1'b0;
    n8007[913] = 1'b0;
    n8007[912] = 1'b0;
    n8007[911] = 1'b0;
    n8007[910] = 1'b0;
    n8007[909] = 1'b0;
    n8007[908] = 1'b0;
    n8007[907] = 1'b0;
    n8007[906] = 1'b0;
    n8007[905] = 1'b0;
    n8007[904] = 1'b0;
    n8007[903] = 1'b0;
    n8007[902] = 1'b0;
    n8007[901] = 1'b0;
    n8007[900] = 1'b0;
    n8007[899] = 1'b0;
    n8007[898] = 1'b0;
    n8007[897] = 1'b0;
    n8007[896] = 1'b0;
    n8007[895] = 1'b0;
    n8007[894] = 1'b0;
    n8007[893] = 1'b0;
    n8007[892] = 1'b0;
    n8007[891] = 1'b0;
    n8007[890] = 1'b0;
    n8007[889] = 1'b0;
    n8007[888] = 1'b0;
    n8007[887] = 1'b0;
    n8007[886] = 1'b0;
    n8007[885] = 1'b0;
    n8007[884] = 1'b0;
    n8007[883] = 1'b0;
    n8007[882] = 1'b0;
    n8007[881] = 1'b0;
    n8007[880] = 1'b0;
    n8007[879] = 1'b0;
    n8007[878] = 1'b0;
    n8007[877] = 1'b0;
    n8007[876] = 1'b0;
    n8007[875] = 1'b0;
    n8007[874] = 1'b0;
    n8007[873] = 1'b0;
    n8007[872] = 1'b0;
    n8007[871] = 1'b0;
    n8007[870] = 1'b0;
    n8007[869] = 1'b0;
    n8007[868] = 1'b0;
    n8007[867] = 1'b0;
    n8007[866] = 1'b0;
    n8007[865] = 1'b0;
    n8007[864] = 1'b0;
    n8007[863] = 1'b0;
    n8007[862] = 1'b0;
    n8007[861] = 1'b0;
    n8007[860] = 1'b0;
    n8007[859] = 1'b0;
    n8007[858] = 1'b0;
    n8007[857] = 1'b0;
    n8007[856] = 1'b0;
    n8007[855] = 1'b0;
    n8007[854] = 1'b0;
    n8007[853] = 1'b0;
    n8007[852] = 1'b0;
    n8007[851] = 1'b0;
    n8007[850] = 1'b0;
    n8007[849] = 1'b0;
    n8007[848] = 1'b0;
    n8007[847] = 1'b0;
    n8007[846] = 1'b0;
    n8007[845] = 1'b0;
    n8007[844] = 1'b0;
    n8007[843] = 1'b0;
    n8007[842] = 1'b0;
    n8007[841] = 1'b0;
    n8007[840] = 1'b0;
    n8007[839] = 1'b0;
    n8007[838] = 1'b0;
    n8007[837] = 1'b0;
    n8007[836] = 1'b0;
    n8007[835] = 1'b0;
    n8007[834] = 1'b0;
    n8007[833] = 1'b0;
    n8007[832] = 1'b0;
    n8007[831] = 1'b0;
    n8007[830] = 1'b0;
    n8007[829] = 1'b0;
    n8007[828] = 1'b0;
    n8007[827] = 1'b0;
    n8007[826] = 1'b0;
    n8007[825] = 1'b0;
    n8007[824] = 1'b0;
    n8007[823] = 1'b0;
    n8007[822] = 1'b0;
    n8007[821] = 1'b0;
    n8007[820] = 1'b0;
    n8007[819] = 1'b0;
    n8007[818] = 1'b0;
    n8007[817] = 1'b0;
    n8007[816] = 1'b0;
    n8007[815] = 1'b0;
    n8007[814] = 1'b0;
    n8007[813] = 1'b0;
    n8007[812] = 1'b0;
    n8007[811] = 1'b0;
    n8007[810] = 1'b0;
    n8007[809] = 1'b0;
    n8007[808] = 1'b0;
    n8007[807] = 1'b0;
    n8007[806] = 1'b0;
    n8007[805] = 1'b0;
    n8007[804] = 1'b0;
    n8007[803] = 1'b0;
    n8007[802] = 1'b0;
    n8007[801] = 1'b0;
    n8007[800] = 1'b0;
    n8007[799] = 1'b0;
    n8007[798] = 1'b0;
    n8007[797] = 1'b0;
    n8007[796] = 1'b0;
    n8007[795] = 1'b0;
    n8007[794] = 1'b0;
    n8007[793] = 1'b0;
    n8007[792] = 1'b0;
    n8007[791] = 1'b0;
    n8007[790] = 1'b0;
    n8007[789] = 1'b0;
    n8007[788] = 1'b0;
    n8007[787] = 1'b0;
    n8007[786] = 1'b0;
    n8007[785] = 1'b0;
    n8007[784] = 1'b0;
    n8007[783] = 1'b0;
    n8007[782] = 1'b0;
    n8007[781] = 1'b0;
    n8007[780] = 1'b0;
    n8007[779] = 1'b0;
    n8007[778] = 1'b0;
    n8007[777] = 1'b0;
    n8007[776] = 1'b0;
    n8007[775] = 1'b0;
    n8007[774] = 1'b0;
    n8007[773] = 1'b0;
    n8007[772] = 1'b0;
    n8007[771] = 1'b0;
    n8007[770] = 1'b0;
    n8007[769] = 1'b0;
    n8007[768] = 1'b0;
    n8007[767] = 1'b0;
    n8007[766] = 1'b0;
    n8007[765] = 1'b0;
    n8007[764] = 1'b0;
    n8007[763] = 1'b0;
    n8007[762] = 1'b0;
    n8007[761] = 1'b0;
    n8007[760] = 1'b0;
    n8007[759] = 1'b0;
    n8007[758] = 1'b0;
    n8007[757] = 1'b0;
    n8007[756] = 1'b0;
    n8007[755] = 1'b0;
    n8007[754] = 1'b0;
    n8007[753] = 1'b0;
    n8007[752] = 1'b0;
    n8007[751] = 1'b0;
    n8007[750] = 1'b0;
    n8007[749] = 1'b0;
    n8007[748] = 1'b0;
    n8007[747] = 1'b0;
    n8007[746] = 1'b0;
    n8007[745] = 1'b0;
    n8007[744] = 1'b0;
    n8007[743] = 1'b0;
    n8007[742] = 1'b0;
    n8007[741] = 1'b0;
    n8007[740] = 1'b0;
    n8007[739] = 1'b0;
    n8007[738] = 1'b0;
    n8007[737] = 1'b0;
    n8007[736] = 1'b0;
    n8007[735] = 1'b0;
    n8007[734] = 1'b0;
    n8007[733] = 1'b0;
    n8007[732] = 1'b0;
    n8007[731] = 1'b0;
    n8007[730] = 1'b0;
    n8007[729] = 1'b0;
    n8007[728] = 1'b0;
    n8007[727] = 1'b0;
    n8007[726] = 1'b0;
    n8007[725] = 1'b0;
    n8007[724] = 1'b0;
    n8007[723] = 1'b0;
    n8007[722] = 1'b0;
    n8007[721] = 1'b0;
    n8007[720] = 1'b0;
    n8007[719] = 1'b0;
    n8007[718] = 1'b0;
    n8007[717] = 1'b0;
    n8007[716] = 1'b0;
    n8007[715] = 1'b0;
    n8007[714] = 1'b0;
    n8007[713] = 1'b0;
    n8007[712] = 1'b0;
    n8007[711] = 1'b0;
    n8007[710] = 1'b0;
    n8007[709] = 1'b0;
    n8007[708] = 1'b0;
    n8007[707] = 1'b0;
    n8007[706] = 1'b0;
    n8007[705] = 1'b0;
    n8007[704] = 1'b0;
    n8007[703] = 1'b0;
    n8007[702] = 1'b0;
    n8007[701] = 1'b0;
    n8007[700] = 1'b0;
    n8007[699] = 1'b0;
    n8007[698] = 1'b0;
    n8007[697] = 1'b0;
    n8007[696] = 1'b0;
    n8007[695] = 1'b0;
    n8007[694] = 1'b0;
    n8007[693] = 1'b0;
    n8007[692] = 1'b0;
    n8007[691] = 1'b0;
    n8007[690] = 1'b0;
    n8007[689] = 1'b0;
    n8007[688] = 1'b0;
    n8007[687] = 1'b0;
    n8007[686] = 1'b0;
    n8007[685] = 1'b0;
    n8007[684] = 1'b0;
    n8007[683] = 1'b0;
    n8007[682] = 1'b0;
    n8007[681] = 1'b0;
    n8007[680] = 1'b0;
    n8007[679] = 1'b0;
    n8007[678] = 1'b0;
    n8007[677] = 1'b0;
    n8007[676] = 1'b0;
    n8007[675] = 1'b0;
    n8007[674] = 1'b0;
    n8007[673] = 1'b0;
    n8007[672] = 1'b0;
    n8007[671] = 1'b0;
    n8007[670] = 1'b0;
    n8007[669] = 1'b0;
    n8007[668] = 1'b0;
    n8007[667] = 1'b0;
    n8007[666] = 1'b0;
    n8007[665] = 1'b0;
    n8007[664] = 1'b0;
    n8007[663] = 1'b0;
    n8007[662] = 1'b0;
    n8007[661] = 1'b0;
    n8007[660] = 1'b0;
    n8007[659] = 1'b0;
    n8007[658] = 1'b0;
    n8007[657] = 1'b0;
    n8007[656] = 1'b0;
    n8007[655] = 1'b0;
    n8007[654] = 1'b0;
    n8007[653] = 1'b0;
    n8007[652] = 1'b0;
    n8007[651] = 1'b0;
    n8007[650] = 1'b0;
    n8007[649] = 1'b0;
    n8007[648] = 1'b0;
    n8007[647] = 1'b0;
    n8007[646] = 1'b0;
    n8007[645] = 1'b0;
    n8007[644] = 1'b0;
    n8007[643] = 1'b0;
    n8007[642] = 1'b0;
    n8007[641] = 1'b0;
    n8007[640] = 1'b0;
    n8007[639] = 1'b0;
    n8007[638] = 1'b0;
    n8007[637] = 1'b0;
    n8007[636] = 1'b0;
    n8007[635] = 1'b0;
    n8007[634] = 1'b0;
    n8007[633] = 1'b0;
    n8007[632] = 1'b0;
    n8007[631] = 1'b0;
    n8007[630] = 1'b0;
    n8007[629] = 1'b0;
    n8007[628] = 1'b0;
    n8007[627] = 1'b0;
    n8007[626] = 1'b0;
    n8007[625] = 1'b0;
    n8007[624] = 1'b0;
    n8007[623] = 1'b0;
    n8007[622] = 1'b0;
    n8007[621] = 1'b0;
    n8007[620] = 1'b0;
    n8007[619] = 1'b0;
    n8007[618] = 1'b0;
    n8007[617] = 1'b0;
    n8007[616] = 1'b0;
    n8007[615] = 1'b0;
    n8007[614] = 1'b0;
    n8007[613] = 1'b0;
    n8007[612] = 1'b0;
    n8007[611] = 1'b0;
    n8007[610] = 1'b0;
    n8007[609] = 1'b0;
    n8007[608] = 1'b0;
    n8007[607] = 1'b0;
    n8007[606] = 1'b0;
    n8007[605] = 1'b0;
    n8007[604] = 1'b0;
    n8007[603] = 1'b0;
    n8007[602] = 1'b0;
    n8007[601] = 1'b0;
    n8007[600] = 1'b0;
    n8007[599] = 1'b0;
    n8007[598] = 1'b0;
    n8007[597] = 1'b0;
    n8007[596] = 1'b0;
    n8007[595] = 1'b0;
    n8007[594] = 1'b0;
    n8007[593] = 1'b0;
    n8007[592] = 1'b0;
    n8007[591] = 1'b0;
    n8007[590] = 1'b0;
    n8007[589] = 1'b0;
    n8007[588] = 1'b0;
    n8007[587] = 1'b0;
    n8007[586] = 1'b0;
    n8007[585] = 1'b0;
    n8007[584] = 1'b0;
    n8007[583] = 1'b0;
    n8007[582] = 1'b0;
    n8007[581] = 1'b0;
    n8007[580] = 1'b0;
    n8007[579] = 1'b0;
    n8007[578] = 1'b0;
    n8007[577] = 1'b0;
    n8007[576] = 1'b0;
    n8007[575] = 1'b0;
    n8007[574] = 1'b0;
    n8007[573] = 1'b0;
    n8007[572] = 1'b0;
    n8007[571] = 1'b0;
    n8007[570] = 1'b0;
    n8007[569] = 1'b0;
    n8007[568] = 1'b0;
    n8007[567] = 1'b0;
    n8007[566] = 1'b0;
    n8007[565] = 1'b0;
    n8007[564] = 1'b0;
    n8007[563] = 1'b0;
    n8007[562] = 1'b0;
    n8007[561] = 1'b0;
    n8007[560] = 1'b0;
    n8007[559] = 1'b0;
    n8007[558] = 1'b0;
    n8007[557] = 1'b0;
    n8007[556] = 1'b0;
    n8007[555] = 1'b0;
    n8007[554] = 1'b0;
    n8007[553] = 1'b0;
    n8007[552] = 1'b0;
    n8007[551] = 1'b0;
    n8007[550] = 1'b0;
    n8007[549] = 1'b0;
    n8007[548] = 1'b0;
    n8007[547] = 1'b0;
    n8007[546] = 1'b0;
    n8007[545] = 1'b0;
    n8007[544] = 1'b0;
    n8007[543] = 1'b0;
    n8007[542] = 1'b0;
    n8007[541] = 1'b0;
    n8007[540] = 1'b0;
    n8007[539] = 1'b0;
    n8007[538] = 1'b0;
    n8007[537] = 1'b0;
    n8007[536] = 1'b0;
    n8007[535] = 1'b0;
    n8007[534] = 1'b0;
    n8007[533] = 1'b0;
    n8007[532] = 1'b0;
    n8007[531] = 1'b0;
    n8007[530] = 1'b0;
    n8007[529] = 1'b0;
    n8007[528] = 1'b0;
    n8007[527] = 1'b0;
    n8007[526] = 1'b0;
    n8007[525] = 1'b0;
    n8007[524] = 1'b0;
    n8007[523] = 1'b0;
    n8007[522] = 1'b0;
    n8007[521] = 1'b0;
    n8007[520] = 1'b0;
    n8007[519] = 1'b0;
    n8007[518] = 1'b0;
    n8007[517] = 1'b0;
    n8007[516] = 1'b0;
    n8007[515] = 1'b0;
    n8007[514] = 1'b0;
    n8007[513] = 1'b0;
    n8007[512] = 1'b0;
    n8007[511] = 1'b1;
    n8007[510] = 1'b1;
    n8007[509] = 1'b1;
    n8007[508] = 1'b1;
    n8007[507] = 1'b1;
    n8007[506] = 1'b1;
    n8007[505] = 1'b1;
    n8007[504] = 1'b1;
    n8007[503] = 1'b1;
    n8007[502] = 1'b1;
    n8007[501] = 1'b1;
    n8007[500] = 1'b1;
    n8007[499] = 1'b1;
    n8007[498] = 1'b1;
    n8007[497] = 1'b1;
    n8007[496] = 1'b1;
    n8007[495] = 1'b1;
    n8007[494] = 1'b1;
    n8007[493] = 1'b1;
    n8007[492] = 1'b1;
    n8007[491] = 1'b1;
    n8007[490] = 1'b1;
    n8007[489] = 1'b1;
    n8007[488] = 1'b1;
    n8007[487] = 1'b1;
    n8007[486] = 1'b1;
    n8007[485] = 1'b1;
    n8007[484] = 1'b1;
    n8007[483] = 1'b1;
    n8007[482] = 1'b1;
    n8007[481] = 1'b1;
    n8007[480] = 1'b1;
    n8007[479] = 1'b1;
    n8007[478] = 1'b1;
    n8007[477] = 1'b1;
    n8007[476] = 1'b1;
    n8007[475] = 1'b1;
    n8007[474] = 1'b1;
    n8007[473] = 1'b1;
    n8007[472] = 1'b1;
    n8007[471] = 1'b1;
    n8007[470] = 1'b1;
    n8007[469] = 1'b1;
    n8007[468] = 1'b1;
    n8007[467] = 1'b1;
    n8007[466] = 1'b1;
    n8007[465] = 1'b1;
    n8007[464] = 1'b1;
    n8007[463] = 1'b1;
    n8007[462] = 1'b1;
    n8007[461] = 1'b1;
    n8007[460] = 1'b1;
    n8007[459] = 1'b1;
    n8007[458] = 1'b1;
    n8007[457] = 1'b1;
    n8007[456] = 1'b1;
    n8007[455] = 1'b1;
    n8007[454] = 1'b1;
    n8007[453] = 1'b1;
    n8007[452] = 1'b1;
    n8007[451] = 1'b1;
    n8007[450] = 1'b1;
    n8007[449] = 1'b1;
    n8007[448] = 1'b1;
    n8007[447] = 1'b0;
    n8007[446] = 1'b0;
    n8007[445] = 1'b0;
    n8007[444] = 1'b0;
    n8007[443] = 1'b0;
    n8007[442] = 1'b0;
    n8007[441] = 1'b0;
    n8007[440] = 1'b0;
    n8007[439] = 1'b0;
    n8007[438] = 1'b0;
    n8007[437] = 1'b0;
    n8007[436] = 1'b0;
    n8007[435] = 1'b0;
    n8007[434] = 1'b0;
    n8007[433] = 1'b0;
    n8007[432] = 1'b0;
    n8007[431] = 1'b0;
    n8007[430] = 1'b0;
    n8007[429] = 1'b0;
    n8007[428] = 1'b0;
    n8007[427] = 1'b0;
    n8007[426] = 1'b0;
    n8007[425] = 1'b0;
    n8007[424] = 1'b0;
    n8007[423] = 1'b0;
    n8007[422] = 1'b0;
    n8007[421] = 1'b0;
    n8007[420] = 1'b0;
    n8007[419] = 1'b0;
    n8007[418] = 1'b0;
    n8007[417] = 1'b0;
    n8007[416] = 1'b0;
    n8007[415] = 1'b1;
    n8007[414] = 1'b1;
    n8007[413] = 1'b1;
    n8007[412] = 1'b1;
    n8007[411] = 1'b1;
    n8007[410] = 1'b1;
    n8007[409] = 1'b1;
    n8007[408] = 1'b1;
    n8007[407] = 1'b1;
    n8007[406] = 1'b1;
    n8007[405] = 1'b1;
    n8007[404] = 1'b1;
    n8007[403] = 1'b1;
    n8007[402] = 1'b1;
    n8007[401] = 1'b1;
    n8007[400] = 1'b1;
    n8007[399] = 1'b1;
    n8007[398] = 1'b1;
    n8007[397] = 1'b1;
    n8007[396] = 1'b1;
    n8007[395] = 1'b1;
    n8007[394] = 1'b1;
    n8007[393] = 1'b1;
    n8007[392] = 1'b1;
    n8007[391] = 1'b1;
    n8007[390] = 1'b1;
    n8007[389] = 1'b1;
    n8007[388] = 1'b1;
    n8007[387] = 1'b1;
    n8007[386] = 1'b1;
    n8007[385] = 1'b1;
    n8007[384] = 1'b1;
    n8007[383] = 1'b0;
    n8007[382] = 1'b0;
    n8007[381] = 1'b0;
    n8007[380] = 1'b0;
    n8007[379] = 1'b0;
    n8007[378] = 1'b0;
    n8007[377] = 1'b0;
    n8007[376] = 1'b0;
    n8007[375] = 1'b0;
    n8007[374] = 1'b0;
    n8007[373] = 1'b0;
    n8007[372] = 1'b0;
    n8007[371] = 1'b0;
    n8007[370] = 1'b0;
    n8007[369] = 1'b0;
    n8007[368] = 1'b0;
    n8007[367] = 1'b0;
    n8007[366] = 1'b0;
    n8007[365] = 1'b0;
    n8007[364] = 1'b0;
    n8007[363] = 1'b0;
    n8007[362] = 1'b0;
    n8007[361] = 1'b0;
    n8007[360] = 1'b0;
    n8007[359] = 1'b0;
    n8007[358] = 1'b0;
    n8007[357] = 1'b0;
    n8007[356] = 1'b0;
    n8007[355] = 1'b0;
    n8007[354] = 1'b0;
    n8007[353] = 1'b0;
    n8007[352] = 1'b0;
    n8007[351] = 1'b0;
    n8007[350] = 1'b0;
    n8007[349] = 1'b0;
    n8007[348] = 1'b0;
    n8007[347] = 1'b0;
    n8007[346] = 1'b0;
    n8007[345] = 1'b0;
    n8007[344] = 1'b0;
    n8007[343] = 1'b0;
    n8007[342] = 1'b0;
    n8007[341] = 1'b0;
    n8007[340] = 1'b0;
    n8007[339] = 1'b0;
    n8007[338] = 1'b0;
    n8007[337] = 1'b0;
    n8007[336] = 1'b0;
    n8007[335] = 1'b0;
    n8007[334] = 1'b0;
    n8007[333] = 1'b0;
    n8007[332] = 1'b0;
    n8007[331] = 1'b0;
    n8007[330] = 1'b0;
    n8007[329] = 1'b0;
    n8007[328] = 1'b0;
    n8007[327] = 1'b0;
    n8007[326] = 1'b0;
    n8007[325] = 1'b0;
    n8007[324] = 1'b0;
    n8007[323] = 1'b0;
    n8007[322] = 1'b0;
    n8007[321] = 1'b0;
    n8007[320] = 1'b0;
    n8007[319] = 1'b0;
    n8007[318] = 1'b0;
    n8007[317] = 1'b0;
    n8007[316] = 1'b0;
    n8007[315] = 1'b0;
    n8007[314] = 1'b0;
    n8007[313] = 1'b0;
    n8007[312] = 1'b0;
    n8007[311] = 1'b0;
    n8007[310] = 1'b0;
    n8007[309] = 1'b0;
    n8007[308] = 1'b0;
    n8007[307] = 1'b0;
    n8007[306] = 1'b0;
    n8007[305] = 1'b0;
    n8007[304] = 1'b0;
    n8007[303] = 1'b0;
    n8007[302] = 1'b0;
    n8007[301] = 1'b0;
    n8007[300] = 1'b0;
    n8007[299] = 1'b0;
    n8007[298] = 1'b0;
    n8007[297] = 1'b0;
    n8007[296] = 1'b0;
    n8007[295] = 1'b0;
    n8007[294] = 1'b0;
    n8007[293] = 1'b0;
    n8007[292] = 1'b0;
    n8007[291] = 1'b0;
    n8007[290] = 1'b0;
    n8007[289] = 1'b0;
    n8007[288] = 1'b0;
    n8007[287] = 1'b0;
    n8007[286] = 1'b0;
    n8007[285] = 1'b0;
    n8007[284] = 1'b0;
    n8007[283] = 1'b0;
    n8007[282] = 1'b0;
    n8007[281] = 1'b0;
    n8007[280] = 1'b0;
    n8007[279] = 1'b0;
    n8007[278] = 1'b0;
    n8007[277] = 1'b0;
    n8007[276] = 1'b0;
    n8007[275] = 1'b0;
    n8007[274] = 1'b0;
    n8007[273] = 1'b0;
    n8007[272] = 1'b0;
    n8007[271] = 1'b0;
    n8007[270] = 1'b0;
    n8007[269] = 1'b0;
    n8007[268] = 1'b0;
    n8007[267] = 1'b0;
    n8007[266] = 1'b0;
    n8007[265] = 1'b0;
    n8007[264] = 1'b0;
    n8007[263] = 1'b0;
    n8007[262] = 1'b0;
    n8007[261] = 1'b0;
    n8007[260] = 1'b0;
    n8007[259] = 1'b0;
    n8007[258] = 1'b0;
    n8007[257] = 1'b0;
    n8007[256] = 1'b0;
    n8007[255] = 1'b0;
    n8007[254] = 1'b0;
    n8007[253] = 1'b0;
    n8007[252] = 1'b0;
    n8007[251] = 1'b0;
    n8007[250] = 1'b0;
    n8007[249] = 1'b0;
    n8007[248] = 1'b0;
    n8007[247] = 1'b0;
    n8007[246] = 1'b0;
    n8007[245] = 1'b0;
    n8007[244] = 1'b0;
    n8007[243] = 1'b0;
    n8007[242] = 1'b0;
    n8007[241] = 1'b0;
    n8007[240] = 1'b0;
    n8007[239] = 1'b0;
    n8007[238] = 1'b0;
    n8007[237] = 1'b0;
    n8007[236] = 1'b0;
    n8007[235] = 1'b0;
    n8007[234] = 1'b0;
    n8007[233] = 1'b0;
    n8007[232] = 1'b0;
    n8007[231] = 1'b0;
    n8007[230] = 1'b0;
    n8007[229] = 1'b0;
    n8007[228] = 1'b0;
    n8007[227] = 1'b0;
    n8007[226] = 1'b0;
    n8007[225] = 1'b0;
    n8007[224] = 1'b0;
    n8007[223] = 1'b0;
    n8007[222] = 1'b0;
    n8007[221] = 1'b0;
    n8007[220] = 1'b0;
    n8007[219] = 1'b0;
    n8007[218] = 1'b0;
    n8007[217] = 1'b0;
    n8007[216] = 1'b0;
    n8007[215] = 1'b0;
    n8007[214] = 1'b0;
    n8007[213] = 1'b0;
    n8007[212] = 1'b0;
    n8007[211] = 1'b0;
    n8007[210] = 1'b0;
    n8007[209] = 1'b0;
    n8007[208] = 1'b0;
    n8007[207] = 1'b0;
    n8007[206] = 1'b0;
    n8007[205] = 1'b0;
    n8007[204] = 1'b0;
    n8007[203] = 1'b0;
    n8007[202] = 1'b0;
    n8007[201] = 1'b0;
    n8007[200] = 1'b0;
    n8007[199] = 1'b0;
    n8007[198] = 1'b0;
    n8007[197] = 1'b0;
    n8007[196] = 1'b0;
    n8007[195] = 1'b0;
    n8007[194] = 1'b0;
    n8007[193] = 1'b0;
    n8007[192] = 1'b0;
    n8007[191] = 1'b0;
    n8007[190] = 1'b0;
    n8007[189] = 1'b0;
    n8007[188] = 1'b0;
    n8007[187] = 1'b0;
    n8007[186] = 1'b0;
    n8007[185] = 1'b0;
    n8007[184] = 1'b0;
    n8007[183] = 1'b0;
    n8007[182] = 1'b0;
    n8007[181] = 1'b0;
    n8007[180] = 1'b0;
    n8007[179] = 1'b0;
    n8007[178] = 1'b0;
    n8007[177] = 1'b0;
    n8007[176] = 1'b0;
    n8007[175] = 1'b0;
    n8007[174] = 1'b0;
    n8007[173] = 1'b0;
    n8007[172] = 1'b0;
    n8007[171] = 1'b0;
    n8007[170] = 1'b0;
    n8007[169] = 1'b0;
    n8007[168] = 1'b0;
    n8007[167] = 1'b0;
    n8007[166] = 1'b0;
    n8007[165] = 1'b0;
    n8007[164] = 1'b0;
    n8007[163] = 1'b0;
    n8007[162] = 1'b0;
    n8007[161] = 1'b0;
    n8007[160] = 1'b0;
    n8007[159] = 1'b0;
    n8007[158] = 1'b0;
    n8007[157] = 1'b0;
    n8007[156] = 1'b0;
    n8007[155] = 1'b0;
    n8007[154] = 1'b0;
    n8007[153] = 1'b0;
    n8007[152] = 1'b0;
    n8007[151] = 1'b0;
    n8007[150] = 1'b0;
    n8007[149] = 1'b0;
    n8007[148] = 1'b0;
    n8007[147] = 1'b0;
    n8007[146] = 1'b0;
    n8007[145] = 1'b0;
    n8007[144] = 1'b0;
    n8007[143] = 1'b0;
    n8007[142] = 1'b0;
    n8007[141] = 1'b0;
    n8007[140] = 1'b0;
    n8007[139] = 1'b0;
    n8007[138] = 1'b0;
    n8007[137] = 1'b0;
    n8007[136] = 1'b0;
    n8007[135] = 1'b0;
    n8007[134] = 1'b0;
    n8007[133] = 1'b0;
    n8007[132] = 1'b0;
    n8007[131] = 1'b0;
    n8007[130] = 1'b0;
    n8007[129] = 1'b0;
    n8007[128] = 1'b0;
    n8007[127] = 1'b0;
    n8007[126] = 1'b0;
    n8007[125] = 1'b0;
    n8007[124] = 1'b0;
    n8007[123] = 1'b0;
    n8007[122] = 1'b0;
    n8007[121] = 1'b0;
    n8007[120] = 1'b0;
    n8007[119] = 1'b0;
    n8007[118] = 1'b0;
    n8007[117] = 1'b0;
    n8007[116] = 1'b0;
    n8007[115] = 1'b0;
    n8007[114] = 1'b0;
    n8007[113] = 1'b0;
    n8007[112] = 1'b0;
    n8007[111] = 1'b0;
    n8007[110] = 1'b0;
    n8007[109] = 1'b0;
    n8007[108] = 1'b0;
    n8007[107] = 1'b0;
    n8007[106] = 1'b0;
    n8007[105] = 1'b0;
    n8007[104] = 1'b0;
    n8007[103] = 1'b0;
    n8007[102] = 1'b0;
    n8007[101] = 1'b0;
    n8007[100] = 1'b0;
    n8007[99] = 1'b0;
    n8007[98] = 1'b0;
    n8007[97] = 1'b0;
    n8007[96] = 1'b0;
    n8007[95] = 1'b0;
    n8007[94] = 1'b0;
    n8007[93] = 1'b0;
    n8007[92] = 1'b0;
    n8007[91] = 1'b0;
    n8007[90] = 1'b0;
    n8007[89] = 1'b0;
    n8007[88] = 1'b0;
    n8007[87] = 1'b0;
    n8007[86] = 1'b0;
    n8007[85] = 1'b0;
    n8007[84] = 1'b0;
    n8007[83] = 1'b0;
    n8007[82] = 1'b0;
    n8007[81] = 1'b0;
    n8007[80] = 1'b0;
    n8007[79] = 1'b0;
    n8007[78] = 1'b0;
    n8007[77] = 1'b0;
    n8007[76] = 1'b0;
    n8007[75] = 1'b0;
    n8007[74] = 1'b0;
    n8007[73] = 1'b0;
    n8007[72] = 1'b0;
    n8007[71] = 1'b0;
    n8007[70] = 1'b0;
    n8007[69] = 1'b0;
    n8007[68] = 1'b0;
    n8007[67] = 1'b0;
    n8007[66] = 1'b0;
    n8007[65] = 1'b0;
    n8007[64] = 1'b0;
    n8007[63] = 1'b0;
    n8007[62] = 1'b0;
    n8007[61] = 1'b0;
    n8007[60] = 1'b0;
    n8007[59] = 1'b0;
    n8007[58] = 1'b0;
    n8007[57] = 1'b0;
    n8007[56] = 1'b0;
    n8007[55] = 1'b0;
    n8007[54] = 1'b0;
    n8007[53] = 1'b0;
    n8007[52] = 1'b0;
    n8007[51] = 1'b0;
    n8007[50] = 1'b0;
    n8007[49] = 1'b0;
    n8007[48] = 1'b0;
    n8007[47] = 1'b0;
    n8007[46] = 1'b0;
    n8007[45] = 1'b0;
    n8007[44] = 1'b0;
    n8007[43] = 1'b0;
    n8007[42] = 1'b0;
    n8007[41] = 1'b0;
    n8007[40] = 1'b0;
    n8007[39] = 1'b0;
    n8007[38] = 1'b0;
    n8007[37] = 1'b0;
    n8007[36] = 1'b0;
    n8007[35] = 1'b0;
    n8007[34] = 1'b0;
    n8007[33] = 1'b0;
    n8007[32] = 1'b0;
    n8007[31] = 1'b0;
    n8007[30] = 1'b0;
    n8007[29] = 1'b0;
    n8007[28] = 1'b0;
    n8007[27] = 1'b0;
    n8007[26] = 1'b0;
    n8007[25] = 1'b0;
    n8007[24] = 1'b0;
    n8007[23] = 1'b0;
    n8007[22] = 1'b0;
    n8007[21] = 1'b0;
    n8007[20] = 1'b0;
    n8007[19] = 1'b0;
    n8007[18] = 1'b0;
    n8007[17] = 1'b0;
    n8007[16] = 1'b0;
    n8007[15] = 1'b0;
    n8007[14] = 1'b0;
    n8007[13] = 1'b0;
    n8007[12] = 1'b0;
    n8007[11] = 1'b0;
    n8007[10] = 1'b0;
    n8007[9] = 1'b0;
    n8007[8] = 1'b0;
    n8007[7] = 1'b0;
    n8007[6] = 1'b0;
    n8007[5] = 1'b0;
    n8007[4] = 1'b0;
    n8007[3] = 1'b0;
    n8007[2] = 1'b0;
    n8007[1] = 1'b0;
    n8007[0] = 1'b0;
    end
  assign n8008_data = n8007[n7448_o];
  /* decode1.vhdl:593:50  */
  /* decode1.vhdl:593:49  */
  reg [43:0] n8009[63:0] ; // memory
  initial begin
    n8009[63] = 44'b00000000000000000000000000000000000000000000;
    n8009[62] = 44'b00000000000000000000000000000000000000000000;
    n8009[61] = 44'b00000000000000000000000000000000000000000000;
    n8009[60] = 44'b00000000000000000000000000000000000000000000;
    n8009[59] = 44'b00000000000000000000000000000000000000000000;
    n8009[58] = 44'b00000000000000000000000000000000000000000000;
    n8009[57] = 44'b00000000000000000000000000000000000000000000;
    n8009[56] = 44'b00000000000000000000000000000000000000000000;
    n8009[55] = 44'b00000000000000000000000000000000000000000000;
    n8009[54] = 44'b00000000000000000000000000000000000000000000;
    n8009[53] = 44'b00000000000000000000000000000000000000000000;
    n8009[52] = 44'b00000000000000000000000000000000000000000000;
    n8009[51] = 44'b00000000000000000000000000000000000000000000;
    n8009[50] = 44'b00000000000000000000000000000000000000000000;
    n8009[49] = 44'b00000000000000000000000000000000000000000000;
    n8009[48] = 44'b00000000000000000000000000000000000000000000;
    n8009[47] = 44'b00000000000000000000000000000000000000000000;
    n8009[46] = 44'b00000000000000000000000000000000000000000000;
    n8009[45] = 44'b00000000000000000000000000000000000000000000;
    n8009[44] = 44'b00000000000000000000000000000000000000000000;
    n8009[43] = 44'b00000000000000000000000000000000000000000000;
    n8009[42] = 44'b00000000000000000000000000000000000000000000;
    n8009[41] = 44'b00000000000000000000000000000000000000000000;
    n8009[40] = 44'b00000000000000000000000000000000000000000000;
    n8009[39] = 44'b00000000000000000000000000000000000000000000;
    n8009[38] = 44'b00000000000000000000000000000000000000000000;
    n8009[37] = 44'b00000000000000000000000000000000000000000000;
    n8009[36] = 44'b00000000000000000000000000000000000000000000;
    n8009[35] = 44'b00000000000000000000000000000000000000000000;
    n8009[34] = 44'b00000000000000000000000000000000000000000000;
    n8009[33] = 44'b00000000000000000000000000000000000000000000;
    n8009[32] = 44'b00000000000000000000000000000000000000000000;
    n8009[31] = 44'b00000000000000000000000000000000000000000000;
    n8009[30] = 44'b00000000000000000000000000000000000000000000;
    n8009[29] = 44'b00000000000000000000000000000000000000000000;
    n8009[28] = 44'b00000000000000000000000000000000000000000000;
    n8009[27] = 44'b00000000000000000000000000000000000000000000;
    n8009[26] = 44'b00000000000000000000000000000000000000000000;
    n8009[25] = 44'b00000000000000000000000000000000000000000000;
    n8009[24] = 44'b00000000000000000000000000000000000000000000;
    n8009[23] = 44'b00000000000000000000000000000000000000000000;
    n8009[22] = 44'b00000000000000000000000000000000000000000000;
    n8009[21] = 44'b00000000000000000000000000000000000000000000;
    n8009[20] = 44'b00000000000000000000000000000000000000000000;
    n8009[19] = 44'b00000000000000000000000000000000000000000000;
    n8009[18] = 44'b00000000000000000000000000000000000000000000;
    n8009[17] = 44'b00000000000000000000000000000000000000000000;
    n8009[16] = 44'b00000000000000000000000000000000000000000000;
    n8009[15] = 44'b00000010000000000000000010100001001101010001;
    n8009[14] = 44'b00000000000000000000000010100001001101010001;
    n8009[13] = 44'b00000000000000000000000000000000000000000000;
    n8009[12] = 44'b00000010000000000000000010100001001101001001;
    n8009[11] = 44'b00000000000000000000000000000000000000000000;
    n8009[10] = 44'b00000000000000000000000000000000000000000000;
    n8009[9] = 44'b00000000000000000000000000000000000000000000;
    n8009[8] = 44'b00000000000000000000000000000000000000000000;
    n8009[7] = 44'b00000000000000000000000000000000000000000000;
    n8009[6] = 44'b00000000000000000000000000000000000000000000;
    n8009[5] = 44'b00000000000000000000000000000000000000000000;
    n8009[4] = 44'b00000000000000000000000000000000000000000000;
    n8009[3] = 44'b00000000000000000000000000000000000000000000;
    n8009[2] = 44'b00000000000000000000000000000000000000000000;
    n8009[1] = 44'b00000000000000000000000000000000000000000000;
    n8009[0] = 44'b00000000000000000000000000000000000000000000;
    end
  assign n8010_data = n8009[n7456_o];
  /* decode1.vhdl:594:43  */
  /* decode1.vhdl:594:42  */
  reg [43:0] n8011[1023:0] ; // memory
  initial begin
    n8011[1023] = 44'b00000010000000001101100000000001001001001001;
    n8011[1022] = 44'b00000000000000000000000000000000000000000000;
    n8011[1021] = 44'b00000000000000000000000000000000000000000000;
    n8011[1020] = 44'b00000000000000000000000000000000000000000000;
    n8011[1019] = 44'b00000001000000000000000000000001001111001001;
    n8011[1018] = 44'b00000000000000000000000000000000000000000000;
    n8011[1017] = 44'b00000000000000000000000000000000000000000000;
    n8011[1016] = 44'b00000000000000000000000000000000000000000000;
    n8011[1015] = 44'b00001000000000011101000010000001001000010001;
    n8011[1014] = 44'b00001000000000000000000010000001001101010001;
    n8011[1013] = 44'b00001000000000010000000010000001001000010001;
    n8011[1012] = 44'b00001001000000000000000010000001001101011001;
    n8011[1011] = 44'b00000000000000000000000000000000000000000000;
    n8011[1010] = 44'b00000000000000000000000000000000000000000000;
    n8011[1009] = 44'b00000000000000000000000000000000000000000000;
    n8011[1008] = 44'b00000000000000000000010010000001010011101001;
    n8011[1007] = 44'b00000000000000000000000000000000000000000000;
    n8011[1006] = 44'b00000000000000000000000000000000000000000000;
    n8011[1005] = 44'b00000000000000000000000000000000000000000000;
    n8011[1004] = 44'b00000000000000000000010010000000000100010001;
    n8011[1003] = 44'b00000000100001100000000010000001010011111010;
    n8011[1002] = 44'b00000000000010000000000010000001010011111010;
    n8011[1001] = 44'b00100000000000000000000000000000000011100001;
    n8011[1000] = 44'b00000000000001100000000010000001010011111010;
    n8011[999] = 44'b00001001000000000000000100010001000110101001;
    n8011[998] = 44'b00000000000000000000000000000000000000000000;
    n8011[997] = 44'b00001001000000000000000100010000000001101001;
    n8011[996] = 44'b00001000000000000000000100010001000110101001;
    n8011[995] = 44'b00001000000000000000000100010001000000011001;
    n8011[994] = 44'b00000000000000000000000000000000000000000000;
    n8011[993] = 44'b00100000000000000000000000000000000000001001;
    n8011[992] = 44'b00000000000000000000000000000000000000000000;
    n8011[991] = 44'b00000000000000001101100000000001001001001001;
    n8011[990] = 44'b00000000000000000000000000000000000000000000;
    n8011[989] = 44'b00000000000000000000000000000000000000000000;
    n8011[988] = 44'b00000000000000000000000000000000000000000000;
    n8011[987] = 44'b00000000000000000000000000000000000000000000;
    n8011[986] = 44'b00000000000000000000000000000000000000000000;
    n8011[985] = 44'b00000000000000000000000000000000000000000000;
    n8011[984] = 44'b00000000000000000000000000000000000000000000;
    n8011[983] = 44'b00001000000000001101000010000001001000010001;
    n8011[982] = 44'b00000000000000000000000000000000000000000000;
    n8011[981] = 44'b00000000000000000000000000000000000000000000;
    n8011[980] = 44'b00000000000000000000000000000000000000000000;
    n8011[979] = 44'b00000000000000000000000000000000000000000000;
    n8011[978] = 44'b00000000000000000000000000000000000000000000;
    n8011[977] = 44'b00000000000000000000000000000000000000000000;
    n8011[976] = 44'b00000000000000000000010010000001010011101001;
    n8011[975] = 44'b00000000000000000000000000000000000000000000;
    n8011[974] = 44'b00000000000000000000000000000000000000000000;
    n8011[973] = 44'b00000000000000000000000000000000000000000000;
    n8011[972] = 44'b00000000000000000000000000000000000000000000;
    n8011[971] = 44'b00000000100000100000000010000001010011111010;
    n8011[970] = 44'b11000000010010000000000010000001010011111010;
    n8011[969] = 44'b00100000000000000000000000000000000010001001;
    n8011[968] = 44'b11000000010001100000000010000001010011111010;
    n8011[967] = 44'b00000000000000000000000000000000000000000000;
    n8011[966] = 44'b00000000000000000000000000000000000000000000;
    n8011[965] = 44'b00001000000000000000000100010000000001101001;
    n8011[964] = 44'b00000000000000000000000000000000000000000000;
    n8011[963] = 44'b00001000000000000001000100010001000000011001;
    n8011[962] = 44'b00000000000000000000000000000000000000000000;
    n8011[961] = 44'b00000000000000000000000000000000000000000000;
    n8011[960] = 44'b00000000000000000000000000000000000000000000;
    n8011[959] = 44'b00000000000000000000000000000000000000000000;
    n8011[958] = 44'b00000000000000000000000000000000000000000000;
    n8011[957] = 44'b00000000000000000000000000000000000000000000;
    n8011[956] = 44'b00000000000000000000000000000000000000000000;
    n8011[955] = 44'b00000000000000000000000000000001001111001001;
    n8011[954] = 44'b00000000000000000000000000000000000000000000;
    n8011[953] = 44'b00000000000000000000000000000000000000000000;
    n8011[952] = 44'b00000000000000000000000000000000000000000000;
    n8011[951] = 44'b00000000000000000000000000000000000000000000;
    n8011[950] = 44'b00001010000000000000000010000001001101010001;
    n8011[949] = 44'b00000000000000000000000010000001001111100001;
    n8011[948] = 44'b00001011000000000000000010000001001101011001;
    n8011[947] = 44'b00000000000000000000000000000000000000000000;
    n8011[946] = 44'b00000000000000000000000000000000000000000000;
    n8011[945] = 44'b00000000000000000000000000000000000000000000;
    n8011[944] = 44'b00000000000000000000010010000001010011101001;
    n8011[943] = 44'b00000000000000000000000000000000000000000000;
    n8011[942] = 44'b00000000000000000000000000000000000000000000;
    n8011[941] = 44'b00000000000000000000000000000000000000000000;
    n8011[940] = 44'b00100000000000000000000010000000000100011001;
    n8011[939] = 44'b00000000100010000000000010000001010011111010;
    n8011[938] = 44'b00000000000000000000000000000000000000000000;
    n8011[937] = 44'b00100000000000000000000000000000000010000001;
    n8011[936] = 44'b00000000000000100000000010000001010011111010;
    n8011[935] = 44'b00000000000000000000000000000000000000000000;
    n8011[934] = 44'b00000000000000000000000000000000000000000000;
    n8011[933] = 44'b00000000000000000000000000000000000000000000;
    n8011[932] = 44'b00000000000000000000000000000000000000000000;
    n8011[931] = 44'b00000000000000000000000000000000000000000000;
    n8011[930] = 44'b00000000000000000000000000000000000000000000;
    n8011[929] = 44'b00000000000000000000000000000000000000000000;
    n8011[928] = 44'b00000000000000000000000000000000000000000000;
    n8011[927] = 44'b00000000000000000000000000000000000000000000;
    n8011[926] = 44'b00000000000000000000000000000000000000000000;
    n8011[925] = 44'b00000000000000000000000000000000000000000000;
    n8011[924] = 44'b00000000000000000000000000000000000000000000;
    n8011[923] = 44'b00000000000000000000000000000000000000000000;
    n8011[922] = 44'b00000000000000000000000000000000000000000000;
    n8011[921] = 44'b00000000000000000000000000000000000000000000;
    n8011[920] = 44'b00000000000000000000000000000000000000000000;
    n8011[919] = 44'b00001000000000001101000010000000001000010001;
    n8011[918] = 44'b00000000000000000000000000000000000000000000;
    n8011[917] = 44'b00000000000000000000000000000000000000000000;
    n8011[916] = 44'b00000000000000000000000000000000000000000000;
    n8011[915] = 44'b00000000000000000000000000000000000000000000;
    n8011[914] = 44'b00000000000000000000000000000000000000000000;
    n8011[913] = 44'b00000000000000000000000000000000000000000000;
    n8011[912] = 44'b00000000000000000000010010000001010011101001;
    n8011[911] = 44'b00000000000000000000000000000000000000000000;
    n8011[910] = 44'b00000000000000000000000000000000000000000000;
    n8011[909] = 44'b00000000000000000000000000000000000000000000;
    n8011[908] = 44'b00000000000000000000000000000000000000000000;
    n8011[907] = 44'b00000000100001000000000010000001010011111010;
    n8011[906] = 44'b00000000000000000000000000000000000000000000;
    n8011[905] = 44'b00000000000000000000000000000000000000000000;
    n8011[904] = 44'b11000000010000100000000010000001010011111010;
    n8011[903] = 44'b00000000000000000000000000000000000000000000;
    n8011[902] = 44'b00000000000000000000000000000000000000000000;
    n8011[901] = 44'b00000000000000100000000100010000000101101001;
    n8011[900] = 44'b00000000000000000000000000000000000000000000;
    n8011[899] = 44'b00001000000000000010000100010001000101100001;
    n8011[898] = 44'b00000000000000000000000000000000000000000000;
    n8011[897] = 44'b00000000000000000000000000000000000000000000;
    n8011[896] = 44'b00000000000000000000000000000000000000000000;
    n8011[895] = 44'b00000000000000000000010010000000000110100001;
    n8011[894] = 44'b00000000000000000000000000000000000000000000;
    n8011[893] = 44'b00000000000000000000000000000000000000000000;
    n8011[892] = 44'b00000000000000000000000000000000000000000000;
    n8011[891] = 44'b00000000000000000000000000000000000000000000;
    n8011[890] = 44'b00000000000000000000000000000000000000000000;
    n8011[889] = 44'b00000000000000000000000000000000000000000000;
    n8011[888] = 44'b00000000000000000000000000000000000000000000;
    n8011[887] = 44'b00001000000000010101000010000001001000010001;
    n8011[886] = 44'b00000000000000000000000000000000000000000000;
    n8011[885] = 44'b00001000000000010100000010000001001000010001;
    n8011[884] = 44'b00000000000000000000000000000000000000000000;
    n8011[883] = 44'b00000000000000000000000000000000000000000000;
    n8011[882] = 44'b00000000000000000000000000000000000000000000;
    n8011[881] = 44'b00000000000000000000000000000000000000000000;
    n8011[880] = 44'b00000000000000000000010010000001010011101001;
    n8011[879] = 44'b00000000000000000000100000010000000100110001;
    n8011[878] = 44'b00000000000000000000000000000000000000000000;
    n8011[877] = 44'b00100001000000000000000000010000000100111001;
    n8011[876] = 44'b00000000000000000000000000000000000000000000;
    n8011[875] = 44'b00000000000000000000000000000000000000000000;
    n8011[874] = 44'b00000000000010000000000000010001010100000010;
    n8011[873] = 44'b00000100100001100000000000010001010100000010;
    n8011[872] = 44'b00000000000001100000000000010001010100000010;
    n8011[871] = 44'b00000000000000000000000000000000000000000000;
    n8011[870] = 44'b00000000000000000000000000000000000000000000;
    n8011[869] = 44'b00000000000001100000000100010000000101110001;
    n8011[868] = 44'b00000000000000000000000000000000000000000000;
    n8011[867] = 44'b00000000000000000000000000000000000000000000;
    n8011[866] = 44'b00000000000000000000000000000000000000000000;
    n8011[865] = 44'b00000000000000000000000000000000000000000000;
    n8011[864] = 44'b00000000000000000000000000000000000000000000;
    n8011[863] = 44'b00000000000000000000000000000000000000000000;
    n8011[862] = 44'b00000000000000000000000000000000000000000000;
    n8011[861] = 44'b00000000000000000000000000000000000000000000;
    n8011[860] = 44'b00000000000000000000000000000000000000000000;
    n8011[859] = 44'b00000000000000000000000000000000000000000000;
    n8011[858] = 44'b00000000000000000000000000000000000000000000;
    n8011[857] = 44'b00000000000000000000000000000000000000000000;
    n8011[856] = 44'b00000000000000000000000000000000000000000000;
    n8011[855] = 44'b00000000000000000000000000000000000000000000;
    n8011[854] = 44'b00000000000000000000000000000000000000000000;
    n8011[853] = 44'b00001000000000011000000010000001001000010001;
    n8011[852] = 44'b00000000000000000000000000000000000000000000;
    n8011[851] = 44'b00000000000000000000000000000000000000000000;
    n8011[850] = 44'b00000000000000000000000000000000000000000000;
    n8011[849] = 44'b00000000000000000000000000000000000000000000;
    n8011[848] = 44'b00000000000000000000010010000001010011101001;
    n8011[847] = 44'b00000000000000000000000000000000000000000000;
    n8011[846] = 44'b00000000000000000000000000000000000000000000;
    n8011[845] = 44'b00100000000000000000000000010000000100111001;
    n8011[844] = 44'b00000000000000000000000000000000000000000000;
    n8011[843] = 44'b00000000000000000000000000000000000000000000;
    n8011[842] = 44'b00000000010010000000000100010001010100000010;
    n8011[841] = 44'b01000100100010000000000000010001010100000010;
    n8011[840] = 44'b00000000010001100000000100010001010100000010;
    n8011[839] = 44'b00000000000000000000000000000000000000000000;
    n8011[838] = 44'b00000000000000000000000000000000000000000000;
    n8011[837] = 44'b00000000000010000000000100010000000101110001;
    n8011[836] = 44'b00000000000000000000000000000000000000000000;
    n8011[835] = 44'b00000000000000000000000000000000000000000000;
    n8011[834] = 44'b00000000000000000000000000000000000000000000;
    n8011[833] = 44'b00000000000000000000000000000000000000000000;
    n8011[832] = 44'b00000000000000000000000000000000000000000000;
    n8011[831] = 44'b00000000000000000000100000000001001001100001;
    n8011[830] = 44'b00000000000000000000000000000000000000000000;
    n8011[829] = 44'b00000000000000000000000000000000000000000000;
    n8011[828] = 44'b00000000000000000000000000000000000000000000;
    n8011[827] = 44'b00000000000000000000000000000000000000000000;
    n8011[826] = 44'b00000000000000000000000000000000000000000000;
    n8011[825] = 44'b00000000000000000000000000000000000000000000;
    n8011[824] = 44'b00000000000000000000000000000000000000000000;
    n8011[823] = 44'b00001000000000010101000010000000001000010001;
    n8011[822] = 44'b00000000000000000000000000000000000000000000;
    n8011[821] = 44'b00001000000000010100000010000000001000010001;
    n8011[820] = 44'b00000000000000000000000000000000000000000000;
    n8011[819] = 44'b00000000000000000000000000000000000000000000;
    n8011[818] = 44'b00000000000000000000000000000000000000000000;
    n8011[817] = 44'b00000000000000000000000000000000000000000000;
    n8011[816] = 44'b00000000000000000000010010000001010011101001;
    n8011[815] = 44'b00000000000000000000000000000000000000000000;
    n8011[814] = 44'b00000000000000000000000000000000000000000000;
    n8011[813] = 44'b00000000000000000000000000000000000000000000;
    n8011[812] = 44'b00000000000000000000000000000000000000000000;
    n8011[811] = 44'b00000000000000000000000000000000000000000000;
    n8011[810] = 44'b00000000000000000000000000000000000000000000;
    n8011[809] = 44'b00000100100010000000000000010001010100000010;
    n8011[808] = 44'b00000000000000100000000000010001010100000010;
    n8011[807] = 44'b00000000000000000000000000000000000000000000;
    n8011[806] = 44'b00000000000000000000000000000000000000000000;
    n8011[805] = 44'b00000000000000000000000000000000000000000000;
    n8011[804] = 44'b00000000000000000000000000000000000000000000;
    n8011[803] = 44'b00000000000000000000000000000000000000000000;
    n8011[802] = 44'b00000000000000000000000000000000000000000000;
    n8011[801] = 44'b00000000000000000000000000000000000000000000;
    n8011[800] = 44'b00000000000000000000000000000000000000000000;
    n8011[799] = 44'b00000000000000000000100000000001001001011001;
    n8011[798] = 44'b00000000000000000000000000000000000000000000;
    n8011[797] = 44'b00000000000000000000000000000000000000000000;
    n8011[796] = 44'b00000000000000000000000000000000000000000000;
    n8011[795] = 44'b00000000000000000000000000000000000000000000;
    n8011[794] = 44'b00000000000000000000000000000000000000000000;
    n8011[793] = 44'b00000000000000000000000000000000000000000000;
    n8011[792] = 44'b00000000000000000000000000000000000000000000;
    n8011[791] = 44'b00001000000000010101000010001011001000010001;
    n8011[790] = 44'b00001010000000000000000010000001001101001001;
    n8011[789] = 44'b00001000000000010100000010001011001000010001;
    n8011[788] = 44'b00001011000000000000000010000001001101001001;
    n8011[787] = 44'b00000000000000000000000000000000000000000000;
    n8011[786] = 44'b00000000000000000000000000000000000000000000;
    n8011[785] = 44'b00000000000000000000000000000000000000000000;
    n8011[784] = 44'b00000000000000000000010010000001010011101001;
    n8011[783] = 44'b00000000000000000000000000000000000000000000;
    n8011[782] = 44'b00000000000000000000000000000000000000000000;
    n8011[781] = 44'b00000000000000000000000000000000000000000000;
    n8011[780] = 44'b00000000000000000000000000000000000000000000;
    n8011[779] = 44'b00000000000000000000000000000000000000000000;
    n8011[778] = 44'b00000000000000000000000000000000000000000000;
    n8011[777] = 44'b00100000000000000000000000000000000010011001;
    n8011[776] = 44'b00000000010000100000000100010001010100000010;
    n8011[775] = 44'b00000000000000000000000000000000000000000000;
    n8011[774] = 44'b00000000000000000000000000000000000000000000;
    n8011[773] = 44'b00000000000000000000000000000000000000000000;
    n8011[772] = 44'b00000000000000000000000000000000000000000000;
    n8011[771] = 44'b00000000000000000000000100010001000001000001;
    n8011[770] = 44'b00000000000000000000000000000000000000000000;
    n8011[769] = 44'b00000000000000000000000000000000000000000000;
    n8011[768] = 44'b00000000000000000000000000000000000000000000;
    n8011[767] = 44'b00000000000000000000000000000000000000000000;
    n8011[766] = 44'b00000000000000000000000000000000000000000000;
    n8011[765] = 44'b00000000000000000000000000000000000000000000;
    n8011[764] = 44'b00000000000000000000000000000000000000000000;
    n8011[763] = 44'b00000000000000000000000000000000000000000000;
    n8011[762] = 44'b00000000000000000000000000000000000000000000;
    n8011[761] = 44'b00000000000000000000000000000000000000000000;
    n8011[760] = 44'b00000000000000000000000000000000000000000000;
    n8011[759] = 44'b00000000000000000000000000000000000000000000;
    n8011[758] = 44'b00000000000000000000000010000001001100101001;
    n8011[757] = 44'b00001000000000000000000010000001001000010001;
    n8011[756] = 44'b00000001000000000000000010000001001100101001;
    n8011[755] = 44'b00000000000000000000000000000000000000000000;
    n8011[754] = 44'b00000000000000000000000000000000000000000000;
    n8011[753] = 44'b00000000000000000000000000000000000000000000;
    n8011[752] = 44'b00000000000000000000010010000001010011101001;
    n8011[751] = 44'b00000000000000000000000000000000000000000000;
    n8011[750] = 44'b00000000000000000000000000000000000000000000;
    n8011[749] = 44'b00000000000000000000000000010001000111000010;
    n8011[748] = 44'b00000000000000000000000000000000000000000000;
    n8011[747] = 44'b10000000100010000000000010000001010011111010;
    n8011[746] = 44'b00000000000000000000000000000000000000000000;
    n8011[745] = 44'b00100000000000000000000000000000000010010001;
    n8011[744] = 44'b00000000000001000000000010000001010011111010;
    n8011[743] = 44'b00000000000000000000000000000000000000000000;
    n8011[742] = 44'b00000000000000000000000000000000000000000000;
    n8011[741] = 44'b00000000000000000001000100010000000111011001;
    n8011[740] = 44'b00000000000000000000000000000000000000000000;
    n8011[739] = 44'b00001000000000000010000100010001000111010001;
    n8011[738] = 44'b00000000000000000000000000000000000000000000;
    n8011[737] = 44'b00000000000000000000000000000000000000000000;
    n8011[736] = 44'b00000000000000000000000000000000000000000000;
    n8011[735] = 44'b00000000000000000000000000000000000000000000;
    n8011[734] = 44'b00000000000000000000000000000000000000000000;
    n8011[733] = 44'b00000000000000000000000000000000000000000000;
    n8011[732] = 44'b00000000000000000000000000000000000000000000;
    n8011[731] = 44'b00000000000000000000000000000000000000000000;
    n8011[730] = 44'b00000000000000000000000000000000000000000000;
    n8011[729] = 44'b00000000000000000000000000000000000000000000;
    n8011[728] = 44'b00000000000000000000000000000000000000000000;
    n8011[727] = 44'b00000000000000000000000000000000000000000000;
    n8011[726] = 44'b00000000000000000000000000000000000000000000;
    n8011[725] = 44'b00000000000000000000000000000000000000000000;
    n8011[724] = 44'b00000000000000000000000000000000000000000000;
    n8011[723] = 44'b00000000000000000000000000000000000000000000;
    n8011[722] = 44'b00000000000000000000000000000000000000000000;
    n8011[721] = 44'b00000000000000000000000000000000000000000000;
    n8011[720] = 44'b00000000000000000000010010000001010011101001;
    n8011[719] = 44'b00000000000000000000000000000000000000000000;
    n8011[718] = 44'b00000000000000000000000000000000000000000000;
    n8011[717] = 44'b00000000000000000000000000010001000111000010;
    n8011[716] = 44'b00000000000000000000000000000000000000000000;
    n8011[715] = 44'b00000000000000000000000000000000000000000000;
    n8011[714] = 44'b00000000000000000000000000000000000000000000;
    n8011[713] = 44'b00000000000000000000000000000000000000000000;
    n8011[712] = 44'b11000000010001000000000010000001010011111010;
    n8011[711] = 44'b00000000000000000000000000000000000000000000;
    n8011[710] = 44'b00000000000000000000000000000000000000000000;
    n8011[709] = 44'b00000000000000000000000100010000000111011001;
    n8011[708] = 44'b00000000000000000000000000000000000000000000;
    n8011[707] = 44'b00001000000000000000000100010001000111010001;
    n8011[706] = 44'b00000000000000000000000000000000000000000000;
    n8011[705] = 44'b00000000000000000000000000000000000000000000;
    n8011[704] = 44'b00000000000000000000000000000000000000000000;
    n8011[703] = 44'b00000000000000000000000000000000000000000000;
    n8011[702] = 44'b00000000000000000000000000000000000000000000;
    n8011[701] = 44'b00000000000000000000000000000000000000000000;
    n8011[700] = 44'b00000000000000000000000000000000000000000000;
    n8011[699] = 44'b00000000000000000000000000000000000000000000;
    n8011[698] = 44'b00000000000000000000000000000000000000000000;
    n8011[697] = 44'b00000000000000000000000000000000000000000000;
    n8011[696] = 44'b00000000000000000000000000000000000000000000;
    n8011[695] = 44'b00000000000000000000000000000000000000000000;
    n8011[694] = 44'b00000000000000000000000000000000000000000000;
    n8011[693] = 44'b00000000000000000000000000000000000000000000;
    n8011[692] = 44'b00000000000000000000000000000000000000000000;
    n8011[691] = 44'b00000000000000000000000000000000000000000000;
    n8011[690] = 44'b00000000000000000000000000000000000000000000;
    n8011[689] = 44'b00000000000000000000000000000000000000000000;
    n8011[688] = 44'b00000000000000000000010010000001010011101001;
    n8011[687] = 44'b00000000000000000000000000000000000000000000;
    n8011[686] = 44'b00000000000000000000000000000000000000000000;
    n8011[685] = 44'b00000000000000000000000000000000000000000000;
    n8011[684] = 44'b00000000000000000000000010010000011100100001;
    n8011[683] = 44'b00000000000000000000000000000000000000000000;
    n8011[682] = 44'b00000000001001100000000010000001010011111010;
    n8011[681] = 44'b00000000000000000000000000000000000000001001;
    n8011[680] = 44'b00000000001001000000000010000001010011111010;
    n8011[679] = 44'b00000000000000000000000000000000000000000000;
    n8011[678] = 44'b00000000000000000000000000000000000000000000;
    n8011[677] = 44'b00000000000000000000000000000000000000000000;
    n8011[676] = 44'b00000000000000000000000000000000000000000000;
    n8011[675] = 44'b00000000000000000000000000000000000000000000;
    n8011[674] = 44'b00000000000000000000000000000000000000000000;
    n8011[673] = 44'b00000000000000000000000000000000000000000000;
    n8011[672] = 44'b00000000000000000000000000000000000000000000;
    n8011[671] = 44'b00000000000000000000000000000000000000000000;
    n8011[670] = 44'b00000000000000000000000000000000000000000000;
    n8011[669] = 44'b00000000000000000000000000000000000000000000;
    n8011[668] = 44'b00000000000000000000000000000000000000000000;
    n8011[667] = 44'b00000000000000000000000000000000000000000000;
    n8011[666] = 44'b00000000000000000000000000000000000000000000;
    n8011[665] = 44'b00000000000000000000000000000000000000000000;
    n8011[664] = 44'b00000000000000000000000000000000000000000000;
    n8011[663] = 44'b00000000000000000000000000000000000000000000;
    n8011[662] = 44'b00000000000000000000000000000000000000000000;
    n8011[661] = 44'b00000000000000000000000000000000000000000000;
    n8011[660] = 44'b00000000000000000000000000000000000000000000;
    n8011[659] = 44'b00000000000000000000000000000000000000000000;
    n8011[658] = 44'b00000000000000000000000000000000000000000000;
    n8011[657] = 44'b00000000000000000000000000000000000000000000;
    n8011[656] = 44'b00000000000000000000010010000001010011101001;
    n8011[655] = 44'b00000000000000000000000000000000000000000000;
    n8011[654] = 44'b00000000000000000000000000000000000000000000;
    n8011[653] = 44'b00000000000000000000000000000000000000000000;
    n8011[652] = 44'b00000000000000000000000000000000000000000000;
    n8011[651] = 44'b00000000000000000000000000000000000000000000;
    n8011[650] = 44'b11000000011001100000000010000001010011111010;
    n8011[649] = 44'b00000000000000000000000000000000000000001001;
    n8011[648] = 44'b11000000011001000000000010000001010011111010;
    n8011[647] = 44'b00000000000000000000000000000000000000000000;
    n8011[646] = 44'b00000000000000000000000000000000000000000000;
    n8011[645] = 44'b00000000000001100000000100010000000101101001;
    n8011[644] = 44'b00000000000000000000000000000000000000000000;
    n8011[643] = 44'b00000000000000000000000000000000000000000000;
    n8011[642] = 44'b00000000000000000000000000000000000000000000;
    n8011[641] = 44'b00000000000000000000000000000000000000000000;
    n8011[640] = 44'b00000000000000000000000000000000000000000000;
    n8011[639] = 44'b00000000000000000000000000000000000000000000;
    n8011[638] = 44'b00000000000000000000000000000000000000000000;
    n8011[637] = 44'b00000000000000000000000000000000000000000000;
    n8011[636] = 44'b00000000000000000000000000000000000000000000;
    n8011[635] = 44'b00000000000000000000000000000000000000000000;
    n8011[634] = 44'b00000000000000000000000000000000000000000000;
    n8011[633] = 44'b00000000000000000000000000000000000000000000;
    n8011[632] = 44'b00000000000000000000000000000000000000000000;
    n8011[631] = 44'b00000000000000000000000000000000000000000000;
    n8011[630] = 44'b00001000000000000000000010000001001010110001;
    n8011[629] = 44'b00000000000000000000000000000000000000000000;
    n8011[628] = 44'b00001001000000000000000010000001001010110001;
    n8011[627] = 44'b00000000000000000000000000000000000000000000;
    n8011[626] = 44'b00000000000000000000000000000000000000000000;
    n8011[625] = 44'b00000000000000000000000000000000000000000000;
    n8011[624] = 44'b00000000000000000000010010000001010011101001;
    n8011[623] = 44'b00000000000000000000000000000000000000000000;
    n8011[622] = 44'b00000000000000000000000000000000000000000000;
    n8011[621] = 44'b00000000000000000000000000000000000000000000;
    n8011[620] = 44'b00000000000000000000000000000000000000000000;
    n8011[619] = 44'b00000000000000000000000000000000000000000000;
    n8011[618] = 44'b00000000000000000000000000000000000000000000;
    n8011[617] = 44'b00000000000000000000000000000000000000000000;
    n8011[616] = 44'b00000000000001000000000000010001010100000010;
    n8011[615] = 44'b00000000000000000000000000000000000000000000;
    n8011[614] = 44'b00000000000000000000000000000000000000000000;
    n8011[613] = 44'b00000000000000000000000000000000000000000000;
    n8011[612] = 44'b00000000000000000000000000000000000000000000;
    n8011[611] = 44'b00001000000000000001000100010001000101100001;
    n8011[610] = 44'b00000000000000000000000000000000000000000000;
    n8011[609] = 44'b00000000000000000000000000000000000000000000;
    n8011[608] = 44'b00000000000000000000000000000000000000000000;
    n8011[607] = 44'b00000000000000000000000000000000000000000000;
    n8011[606] = 44'b00000000000000000000000000000000000000000000;
    n8011[605] = 44'b00000000000000000000000000000000000000000000;
    n8011[604] = 44'b00000000000000000000000000000000000000000000;
    n8011[603] = 44'b00000000000000000000000000000000000000000000;
    n8011[602] = 44'b00000000000000000000000000000000000000000000;
    n8011[601] = 44'b00000000000000000000000000000000000000000000;
    n8011[600] = 44'b00000000000000000000000000000000000000000000;
    n8011[599] = 44'b00000000000000000000000000000000000000000000;
    n8011[598] = 44'b00001010000000000000000010000001001010110001;
    n8011[597] = 44'b00000000000000000000000000000000000000000000;
    n8011[596] = 44'b00001011000000000000000010000001001010110001;
    n8011[595] = 44'b00000000000000000000000000000000000000000000;
    n8011[594] = 44'b00000000000000000000000000000000000000000000;
    n8011[593] = 44'b00000000000000000000000000000000000000000000;
    n8011[592] = 44'b00000000000000000000010010000001010011101001;
    n8011[591] = 44'b00000000000000000000000000000000000000000000;
    n8011[590] = 44'b00000000000000000000000000000000000000000000;
    n8011[589] = 44'b00000000000000000000000000000000000000000000;
    n8011[588] = 44'b00000000000000000000000000000000000000000000;
    n8011[587] = 44'b00000000000000000000000000000000000000000000;
    n8011[586] = 44'b00000000000000000000000000000000000000000000;
    n8011[585] = 44'b00000000000000000000000000000000000000000000;
    n8011[584] = 44'b00000000010001000000000100010001010100000010;
    n8011[583] = 44'b00000000000000000000000000000000000000000000;
    n8011[582] = 44'b00000000000000000000000000000000000000000000;
    n8011[581] = 44'b00000000000000000000000000000000000000000000;
    n8011[580] = 44'b00000000000000000000000000000000000000000000;
    n8011[579] = 44'b00001000000000000000000100010001000101100001;
    n8011[578] = 44'b00000000000000000000000000000000000000000000;
    n8011[577] = 44'b00000000000000000000000000000000000000000000;
    n8011[576] = 44'b00000000000000000000000000000000000000000000;
    n8011[575] = 44'b00000000000000000000000000000000000000000000;
    n8011[574] = 44'b00000000000000000000000000000000000000000000;
    n8011[573] = 44'b00000000000000000000000000000000000000000000;
    n8011[572] = 44'b00000000000000000000000000000000000000000000;
    n8011[571] = 44'b00000000000000000000000000000000000000000000;
    n8011[570] = 44'b00000000000000000000000000000000000000000000;
    n8011[569] = 44'b00000000000000000000000000000000000000000000;
    n8011[568] = 44'b00000000000000000000000000000000000000000000;
    n8011[567] = 44'b00000000000000000000000000000000000000000000;
    n8011[566] = 44'b00001000000000000000000010000001001010101001;
    n8011[565] = 44'b00000000000000000000000000000000000000000000;
    n8011[564] = 44'b00001001000000000000000010000001001010101001;
    n8011[563] = 44'b00000000000000000000000000000000000000000000;
    n8011[562] = 44'b00000000000000000000000000000000000000000000;
    n8011[561] = 44'b00000000000000000000000000000000000000000000;
    n8011[560] = 44'b00000000000000000000010010000001010011101001;
    n8011[559] = 44'b00000000000000000000000000000000000000000000;
    n8011[558] = 44'b00000000000000000000000000000000000000000000;
    n8011[557] = 44'b00000000000000000000000000000000000000000000;
    n8011[556] = 44'b00000000000000000000000110010000000101000001;
    n8011[555] = 44'b00000000000000000000000000000000000000000000;
    n8011[554] = 44'b00000000000000000000000000000000000000000000;
    n8011[553] = 44'b00000000000000000000000000000000000000000000;
    n8011[552] = 44'b00000000000000000000000000000000000000000000;
    n8011[551] = 44'b00000000000000000000000000000000000000000000;
    n8011[550] = 44'b00000000000000000000000000000000000000000000;
    n8011[549] = 44'b00000000000000000000000000000000000000000000;
    n8011[548] = 44'b00000000000000000000000000000000000000000000;
    n8011[547] = 44'b00001000000000000010000100010001000000011001;
    n8011[546] = 44'b00000000000000000000000000000000000000000000;
    n8011[545] = 44'b00000000000000000000000000000000000000000000;
    n8011[544] = 44'b00000000000000000000000000000000000000000000;
    n8011[543] = 44'b00000000000000000000000000000000000000000000;
    n8011[542] = 44'b00000000000000000000000000000000000000000000;
    n8011[541] = 44'b00000000000000000000000000000000000000000000;
    n8011[540] = 44'b00000000000000000000000000000000000000000000;
    n8011[539] = 44'b00000000000000000000000000000000000000000000;
    n8011[538] = 44'b00000000000000000000000000000000000000000000;
    n8011[537] = 44'b00000000000000000000000000000000000000000000;
    n8011[536] = 44'b00000000000000000000000000000000000000000000;
    n8011[535] = 44'b00000000000000000000000000000000000000000000;
    n8011[534] = 44'b00001010000000000000000010000001001010101001;
    n8011[533] = 44'b00000000000000000000000000000000000000000000;
    n8011[532] = 44'b00001011000000000000000010000001001010101001;
    n8011[531] = 44'b00000000000000000000000000000000000000000000;
    n8011[530] = 44'b00000000000000000000000000000000000000000000;
    n8011[529] = 44'b00000000000000000000000000000000000000000000;
    n8011[528] = 44'b00000000000000000000010010000001010011101001;
    n8011[527] = 44'b00000000000000000000000000000000000000000000;
    n8011[526] = 44'b00000000000000000000000000000000000000000000;
    n8011[525] = 44'b00000000000000000000000000000000000111000010;
    n8011[524] = 44'b00000000000000000000000000000000000000000000;
    n8011[523] = 44'b00000000000000000000000000000000000000000000;
    n8011[522] = 44'b00000000000000000000000000000000000000000000;
    n8011[521] = 44'b00000000000000000000000000000000000000000000;
    n8011[520] = 44'b00000000000000000000000000000000000000000000;
    n8011[519] = 44'b00000000000000000000000000000000000000000000;
    n8011[518] = 44'b00000000000000000000000000000000000000000000;
    n8011[517] = 44'b00000000000010000000000100010000000101101001;
    n8011[516] = 44'b00000000000000000000000000000000000000000000;
    n8011[515] = 44'b00000000000000000000000100010001000001010001;
    n8011[514] = 44'b00000000000000000000000000000000000000000000;
    n8011[513] = 44'b00000000000000000000000000000000000000000000;
    n8011[512] = 44'b00000000000000000000000000000000000000000000;
    n8011[511] = 44'b00000000000000000000000000000000000000000000;
    n8011[510] = 44'b00000000000000000000000000000000000000000000;
    n8011[509] = 44'b00000000000000000000000000000000000000000000;
    n8011[508] = 44'b00000000000000000000000000000000000000000000;
    n8011[507] = 44'b00000000000000000000000000000000000000000000;
    n8011[506] = 44'b00000000000000000000000000000000000000000000;
    n8011[505] = 44'b00000000000000000000000000000000000000000000;
    n8011[504] = 44'b00000000000000000000000000000000000000000000;
    n8011[503] = 44'b00001000000000011101000010000001001000010001;
    n8011[502] = 44'b00001000000000000000000010000001001101010001;
    n8011[501] = 44'b00001000000000010000000010000001001000010001;
    n8011[500] = 44'b00001001000000000000000010000001001101011001;
    n8011[499] = 44'b00000000000000000000000000000000000000000000;
    n8011[498] = 44'b00000000000000000000000000000000000000000000;
    n8011[497] = 44'b00000000000000000000000000000000000000000000;
    n8011[496] = 44'b00000000000000000000010010000001010011101001;
    n8011[495] = 44'b00000000000000000000000000000000000000000000;
    n8011[494] = 44'b00000000000000000000000000000000000000000000;
    n8011[493] = 44'b00000000000000000000000000000000000000001001;
    n8011[492] = 44'b00000000000000000000000000000000000000000000;
    n8011[491] = 44'b00000000000110000000000010000001010011111010;
    n8011[490] = 44'b00000000000000000000000000000000000000000000;
    n8011[489] = 44'b00000000000101100000000010000001010011111010;
    n8011[488] = 44'b00000001000001100000001000000001010011111110;
    n8011[487] = 44'b00001001000000000000000100010001000110110001;
    n8011[486] = 44'b00000000000000000000000000000000000000000000;
    n8011[485] = 44'b00001001000000000000000100010000000001101001;
    n8011[484] = 44'b00001000000000000000000100010001000110110001;
    n8011[483] = 44'b00000000000000000000000000000000000000000000;
    n8011[482] = 44'b00000000000000000000000000000000000000000000;
    n8011[481] = 44'b00000000000000000000000000000000000000000000;
    n8011[480] = 44'b00000000000000000000000000000000000000000000;
    n8011[479] = 44'b00000000000000000000000000000000000000000000;
    n8011[478] = 44'b00000000000000000000000000000000000000000000;
    n8011[477] = 44'b00000000000000000000000000000000000000000000;
    n8011[476] = 44'b00000000000000000000000000000000000000000000;
    n8011[475] = 44'b00000000000000000000000000000000000000000000;
    n8011[474] = 44'b00000000000000000000000000000000000000000000;
    n8011[473] = 44'b00000000000000000000000000000000000000000000;
    n8011[472] = 44'b00000000000000000000000000000000000000000000;
    n8011[471] = 44'b00001000000000001101000010000001001000010001;
    n8011[470] = 44'b00000000000000000000000000000000000000000000;
    n8011[469] = 44'b00000000000000000000000000000000000000000000;
    n8011[468] = 44'b00000000000000000000000000000000000000000000;
    n8011[467] = 44'b00000000000000000000000000000000000000000000;
    n8011[466] = 44'b00000000000000000000000000000000000000000000;
    n8011[465] = 44'b00000000000000000000000000000000000000000000;
    n8011[464] = 44'b00000000000000000000010010000001010011101001;
    n8011[463] = 44'b00000000000000000000000000000000000000000000;
    n8011[462] = 44'b00000000000000000000000000000000000000000000;
    n8011[461] = 44'b00000000000000000000000000000000000000001001;
    n8011[460] = 44'b00000000000000000000000000000000000000000000;
    n8011[459] = 44'b00000000000000000000000000000000000000000000;
    n8011[458] = 44'b00000000000000000000000000000000000000000000;
    n8011[457] = 44'b00100000000000000000000000000000000000001001;
    n8011[456] = 44'b11000001010001100000001000000001010011111110;
    n8011[455] = 44'b00000000000000000000000000000000000000000000;
    n8011[454] = 44'b00000000000000000000000000000000000000000000;
    n8011[453] = 44'b00001000000000000000000100010000000001101001;
    n8011[452] = 44'b00000000000000000000000000000000000000000000;
    n8011[451] = 44'b00000000000000000000000000000000000000000000;
    n8011[450] = 44'b00000000000000000000000000000000000000000000;
    n8011[449] = 44'b00000000000000000000000000000000000000000000;
    n8011[448] = 44'b00000000000000000000000000000000000000000000;
    n8011[447] = 44'b00000000000000000000100000000000000100001001;
    n8011[446] = 44'b00000000000000000000000000000000000000000000;
    n8011[445] = 44'b00000000000000000000000000000000000000000000;
    n8011[444] = 44'b00000000000000000000000000000000000000000000;
    n8011[443] = 44'b00000000000000000000000000000000000000000000;
    n8011[442] = 44'b00000000000000000000000000000000000000000000;
    n8011[441] = 44'b00000000000000000000000000000000000000000000;
    n8011[440] = 44'b00000000000000000000000000000000000000000000;
    n8011[439] = 44'b00000000000000000000000000000000000000000000;
    n8011[438] = 44'b00001010000000000000000010000001001101010001;
    n8011[437] = 44'b00000000000000000000000000000000000000000000;
    n8011[436] = 44'b00001011000000000000000010000001001101011001;
    n8011[435] = 44'b00000000000000000000000000000000000000000000;
    n8011[434] = 44'b00000000000000000000000000000000000000000000;
    n8011[433] = 44'b00000000000000000000000000000000000000000000;
    n8011[432] = 44'b00000000000000000000010010000001010011101001;
    n8011[431] = 44'b00000000000000000000000000000000000000000000;
    n8011[430] = 44'b00000000000000000000000000000000000000000000;
    n8011[429] = 44'b00000000000000000000000000000000000000001001;
    n8011[428] = 44'b00000000000000000000000000000000000000000000;
    n8011[427] = 44'b00000000000000000000000000000000000000000000;
    n8011[426] = 44'b00000000000000000000000000000000000000000000;
    n8011[425] = 44'b00100000000000000000000000000000000000001001;
    n8011[424] = 44'b00000000000010000000001000000001010011111110;
    n8011[423] = 44'b00000000000000000000000000000000000000000000;
    n8011[422] = 44'b00000000000000000000000000000000000000000000;
    n8011[421] = 44'b00000000000000000000000000000000000000000000;
    n8011[420] = 44'b00000000000000000000000000000000000000000000;
    n8011[419] = 44'b00000000000000000000000000000000000000000000;
    n8011[418] = 44'b00000000000000000000000000000000000000000000;
    n8011[417] = 44'b00000000000000000000000000000000000000000000;
    n8011[416] = 44'b00000000000000000000000000000000000000000000;
    n8011[415] = 44'b00000000000000000000000000000000000000000000;
    n8011[414] = 44'b00000000000000000000000000000000000000000000;
    n8011[413] = 44'b00000000000000000000000000000000000000000000;
    n8011[412] = 44'b00000000000000000000000000000000000000000000;
    n8011[411] = 44'b00000000000000000000000000000000000000000000;
    n8011[410] = 44'b00000000000000000000000000000000000000000000;
    n8011[409] = 44'b00000000000000000000000000000000000000000000;
    n8011[408] = 44'b00000000000000000000000000000000000000000000;
    n8011[407] = 44'b00001000000000001101000010000000001000010001;
    n8011[406] = 44'b00000000000000000000000000000000000000000000;
    n8011[405] = 44'b00000000000000000000000000000000000000000000;
    n8011[404] = 44'b00000000000000000000000000000000000000000000;
    n8011[403] = 44'b00000000000000000000000000000000000000000000;
    n8011[402] = 44'b00000000000000000000000000000000000000000000;
    n8011[401] = 44'b00000000000000000000000000000000000000000000;
    n8011[400] = 44'b00000000000000000000010010000001010011101001;
    n8011[399] = 44'b00000000000000000000000000000000000000000000;
    n8011[398] = 44'b00000000000000000000000000000000000000000000;
    n8011[397] = 44'b00000000000000000000000000000000000000001001;
    n8011[396] = 44'b00000000000000000000000000000000000000000000;
    n8011[395] = 44'b00000000000000000000000000000000000000000000;
    n8011[394] = 44'b00000000000000000000000000000000000000000000;
    n8011[393] = 44'b00000000000000000000000000000000000000000000;
    n8011[392] = 44'b11000000010010000000001000000001010011111110;
    n8011[391] = 44'b00000000000000000000000000000000000000000000;
    n8011[390] = 44'b00000000000000000000000000000000000000000000;
    n8011[389] = 44'b00000000000000000000000000000000000000000000;
    n8011[388] = 44'b00000000000000000000000000000000000000000000;
    n8011[387] = 44'b00000000000000000000000000000000000000000000;
    n8011[386] = 44'b00000000000000000000000000000000000000000000;
    n8011[385] = 44'b00000000000000000000000000000000000000000000;
    n8011[384] = 44'b00000000000000000000000000000000000000000000;
    n8011[383] = 44'b00000000000000000000000000000000000000000000;
    n8011[382] = 44'b00000000000000000000000000000000000000000000;
    n8011[381] = 44'b00000000000000000000000000000000000000000000;
    n8011[380] = 44'b00000000000000000000000000000000000000000000;
    n8011[379] = 44'b00000000000000000000000000000000000000000000;
    n8011[378] = 44'b00000000000000000000000000000000000000000000;
    n8011[377] = 44'b00000000000000000000000000000000000000000000;
    n8011[376] = 44'b00000000000000000000000000000000000000000000;
    n8011[375] = 44'b00001000000000010101000010000001001000010001;
    n8011[374] = 44'b00000000000000000000000000000000000000000000;
    n8011[373] = 44'b00001000000000010100000010000001001000010001;
    n8011[372] = 44'b00000000000000000000000000000000000000000000;
    n8011[371] = 44'b00000000000000000000000000000000000000000000;
    n8011[370] = 44'b00000000000000000000000000000000000000000000;
    n8011[369] = 44'b00000000000000000000000000000000000000000000;
    n8011[368] = 44'b00000000000000000000010010000001010011101001;
    n8011[367] = 44'b00000000000000000000000000000000000000000000;
    n8011[366] = 44'b00000000000000000000000000000000000000000000;
    n8011[365] = 44'b00000000000000000000000000000000000000001001;
    n8011[364] = 44'b00000000000000000000000000000000000000000000;
    n8011[363] = 44'b00000000000110000000000000010001010100000010;
    n8011[362] = 44'b00000000000000000000000000000000000000000000;
    n8011[361] = 44'b00000000000101100000000000010001010100000010;
    n8011[360] = 44'b00000001000001100000000001000001010100000110;
    n8011[359] = 44'b00000000000000000000000000000000000000000000;
    n8011[358] = 44'b00000000000000000000000000000000000000000000;
    n8011[357] = 44'b00000000000000000000000000000000000000000000;
    n8011[356] = 44'b00000000000000000000000000000000000000000000;
    n8011[355] = 44'b00000000000000000000000000000000000000000000;
    n8011[354] = 44'b00000000000000000000000000000000000000000000;
    n8011[353] = 44'b00000000000000000000000000000000000000000000;
    n8011[352] = 44'b00000000000000000000000000000000000000000000;
    n8011[351] = 44'b00000000000000000000000000000000000000000000;
    n8011[350] = 44'b00000000000000000000000000000000000000000000;
    n8011[349] = 44'b00000000000000000000000000000000000000000000;
    n8011[348] = 44'b00000000000000000000000000000000000000000000;
    n8011[347] = 44'b00000000000000000000000000000000000000000000;
    n8011[346] = 44'b00000000000000000000000000000000000000000000;
    n8011[345] = 44'b00000000000000000000000000000000000000000000;
    n8011[344] = 44'b00000000000000000000000000000000000000000000;
    n8011[343] = 44'b00000000000000000000000000000000000000000000;
    n8011[342] = 44'b00000000000000000000000000000000000000000000;
    n8011[341] = 44'b00000000000000000000000000000000000000000000;
    n8011[340] = 44'b00000000000000000000000000000000000000000000;
    n8011[339] = 44'b00000000000000000000000000000000000000000000;
    n8011[338] = 44'b00000000000000000000000000000000000000000000;
    n8011[337] = 44'b00000000000000000000000000000000000000000000;
    n8011[336] = 44'b00000000000000000000010010000001010011101001;
    n8011[335] = 44'b00000000000000000000000000000000000000000000;
    n8011[334] = 44'b00000000000000000000000000000000000000000000;
    n8011[333] = 44'b00000000000000000000000000000000000000001001;
    n8011[332] = 44'b00000000000000000000000000000000000000000000;
    n8011[331] = 44'b00000000000000000000000000000000000000000000;
    n8011[330] = 44'b00000000000000000000000000000000000000000000;
    n8011[329] = 44'b00000100100000100000000000010001010100000010;
    n8011[328] = 44'b00000001010001100000000101000001010100000110;
    n8011[327] = 44'b00000000000000000000000000000000000000000000;
    n8011[326] = 44'b00000000000000000000000000000000000000000000;
    n8011[325] = 44'b00000000000000000000000000000000000000000000;
    n8011[324] = 44'b00000000000000000000000000000000000000000000;
    n8011[323] = 44'b00000000000000000000000000000000000000000000;
    n8011[322] = 44'b00000000000000000000000000000000000000000000;
    n8011[321] = 44'b00000000000000000000000000000000000000000000;
    n8011[320] = 44'b00000000000000000000000000000000000000000000;
    n8011[319] = 44'b00000000000000000000000000000000000000000000;
    n8011[318] = 44'b00000000000000000000000000000000000000000000;
    n8011[317] = 44'b00000000000000000000000000000000000000000000;
    n8011[316] = 44'b00000000000000000000000000000000000000000000;
    n8011[315] = 44'b00000000000000000000000000000000000000000000;
    n8011[314] = 44'b00000000000000000000000000000000000000000000;
    n8011[313] = 44'b00000000000000000000000000000000000000000000;
    n8011[312] = 44'b00000000000000000000000000000000000000000000;
    n8011[311] = 44'b00001000000000010101000010000000001000010001;
    n8011[310] = 44'b00000000000000000000000000000000000000000000;
    n8011[309] = 44'b00001000000000010100000010000000001000010001;
    n8011[308] = 44'b00000000000000000000000000000000000000000000;
    n8011[307] = 44'b00000000000000000000000000000000000000000000;
    n8011[306] = 44'b00000000000000000000000000000000000000000000;
    n8011[305] = 44'b00000000000000000000000000000000000000000000;
    n8011[304] = 44'b00000000000000000000010010000001010011101001;
    n8011[303] = 44'b00000000000000000000000000000000000000000000;
    n8011[302] = 44'b00000000000000000000000000000000000000000000;
    n8011[301] = 44'b00000000000000000000000000000000000000001001;
    n8011[300] = 44'b00000000000000000000000000000000000000000000;
    n8011[299] = 44'b00000000000000000000000000000000000000000000;
    n8011[298] = 44'b00000000000000000000000000000000000000000000;
    n8011[297] = 44'b00000100100001000000000000010001010100000010;
    n8011[296] = 44'b00000000000010000000000001000001010100000110;
    n8011[295] = 44'b00000000000000000000000000000000000000000000;
    n8011[294] = 44'b00000000000000000000000000000000000000000000;
    n8011[293] = 44'b00000000000000000000000000000000000000000000;
    n8011[292] = 44'b00000000000000000000000000000000000000000000;
    n8011[291] = 44'b00000000000000000000000000000000000000000000;
    n8011[290] = 44'b00000000000000000000000000000000000000000000;
    n8011[289] = 44'b00000000000000000000000000000000000000000000;
    n8011[288] = 44'b00000000000000000000000000000000000000000000;
    n8011[287] = 44'b00000000000000000000000000000000000000000000;
    n8011[286] = 44'b00000000000000000000000000000000000000000000;
    n8011[285] = 44'b00000000000000000000000000000000000000000000;
    n8011[284] = 44'b00000000000000000000000000000000000000000000;
    n8011[283] = 44'b00000000000000000000000000000000000000000000;
    n8011[282] = 44'b00000000000000000000000000000000000000000000;
    n8011[281] = 44'b00000000000000000000000000000000000000000000;
    n8011[280] = 44'b00000000000000000000000000000000000000000000;
    n8011[279] = 44'b00001000000000010101000010001011001000010001;
    n8011[278] = 44'b00001010000000000000000010000001001101001001;
    n8011[277] = 44'b00001000000000010100000010001011001000010001;
    n8011[276] = 44'b00001011000000000000000010000001001101001001;
    n8011[275] = 44'b00000000000000000000000000000000000000000000;
    n8011[274] = 44'b00000000000000000000000000000000000000000000;
    n8011[273] = 44'b00000000000000000000000000000000000000000000;
    n8011[272] = 44'b00000000000000000000010010000001010011101001;
    n8011[271] = 44'b00000000000000000000000000000000000000000000;
    n8011[270] = 44'b00000000000000000000000000000000000000000000;
    n8011[269] = 44'b00000000000000000000000000000000000000001001;
    n8011[268] = 44'b00000000000000000000000010000000000001111001;
    n8011[267] = 44'b00000000000000000000000000000000000000000000;
    n8011[266] = 44'b00000000000000000000000000000000000000000000;
    n8011[265] = 44'b00000000000000000000000000000000000000000000;
    n8011[264] = 44'b00000000010010000000000101000001010100000110;
    n8011[263] = 44'b00000000000000000000000000000000000000000000;
    n8011[262] = 44'b00000000000000000000000000000000000000000000;
    n8011[261] = 44'b00000000000000000000000000000000000000000000;
    n8011[260] = 44'b00000000000000000000000000000000000000000000;
    n8011[259] = 44'b00000000000000000000000000000000000000000000;
    n8011[258] = 44'b00000000000000000000000000000000000000000000;
    n8011[257] = 44'b00000000000000000000000000000000000000000000;
    n8011[256] = 44'b00000000000000000000000000000000000000000000;
    n8011[255] = 44'b00000000000000000000000000000000000000000000;
    n8011[254] = 44'b00000000000000000000000000000000000000000000;
    n8011[253] = 44'b00000000000000000000000000000000000000000000;
    n8011[252] = 44'b00000000000000000000000000000000000000000000;
    n8011[251] = 44'b00000000000000000000000000000000000000000000;
    n8011[250] = 44'b00000000000000000000000000000000000000000000;
    n8011[249] = 44'b00000000000000000000000000000000000000000000;
    n8011[248] = 44'b00000000000000000000000000000000000000000000;
    n8011[247] = 44'b00000000000000000000000000000000000000000000;
    n8011[246] = 44'b00000010000000000000000010000001001100101001;
    n8011[245] = 44'b00001000000000000000000010000001001000010001;
    n8011[244] = 44'b00000011000000000000000010000001001100101001;
    n8011[243] = 44'b00000000000000000000000000000000000000000000;
    n8011[242] = 44'b00000000000000000000000000000000000000000000;
    n8011[241] = 44'b00000000000000000000000000000000000000000000;
    n8011[240] = 44'b00000000000000000000010010000001010011101001;
    n8011[239] = 44'b00000000000000000000000000000000000000000000;
    n8011[238] = 44'b00000000000000000000000000000000000000000000;
    n8011[237] = 44'b00000000000000000000000000000000000000000000;
    n8011[236] = 44'b00000000000000000000000000000000000000000000;
    n8011[235] = 44'b00000000000000000000000000000000000000000000;
    n8011[234] = 44'b00000000000001100000000010000001010011111010;
    n8011[233] = 44'b00000000000101000000000010000001010011111010;
    n8011[232] = 44'b00000000000000000000000000000000000000000000;
    n8011[231] = 44'b00001011000000010000000100010001000110110001;
    n8011[230] = 44'b00000000000000000000000000000000000000000000;
    n8011[229] = 44'b00001010000000010000000100010001000110110001;
    n8011[228] = 44'b00000000000000000000000000000000000000000000;
    n8011[227] = 44'b00000000000000000000000000000000000000000000;
    n8011[226] = 44'b00000000000000000000000000000000000000000000;
    n8011[225] = 44'b00000000000000000000000000000000000000000000;
    n8011[224] = 44'b00000000000000000000000000000000000000000000;
    n8011[223] = 44'b00000000000000000000000000000000000000000000;
    n8011[222] = 44'b00000000000000000000000000000000000000000000;
    n8011[221] = 44'b00000000000000000000000000000000000000000000;
    n8011[220] = 44'b00000000000000000000000000000000000000000000;
    n8011[219] = 44'b00000000000000000000000000000000000000000000;
    n8011[218] = 44'b00000000000000000000000000000000000000000000;
    n8011[217] = 44'b00000000000000000000000000000000000000000000;
    n8011[216] = 44'b00000000000000000000000000000000000000000000;
    n8011[215] = 44'b00000000000000000000000000000000000000000000;
    n8011[214] = 44'b00000000000000000000000000000000000000000000;
    n8011[213] = 44'b00000000000000000000000000000000000000000000;
    n8011[212] = 44'b00000000000000000000000000000000000000000000;
    n8011[211] = 44'b00000000000000000000000000000000000000000000;
    n8011[210] = 44'b00000000000000000000000000000000000000000000;
    n8011[209] = 44'b00000000000000000000000000000000000000000000;
    n8011[208] = 44'b00000000000000000000010010000001010011101001;
    n8011[207] = 44'b00000000000000000000000000000000000000000000;
    n8011[206] = 44'b00000000000000000000000000000000000000000000;
    n8011[205] = 44'b00000000000000000000000000000000000000000000;
    n8011[204] = 44'b00000000000000000000000000000000000000000000;
    n8011[203] = 44'b00000000000000000000000000000000000000000000;
    n8011[202] = 44'b00000000000001000000000010000001010011111010;
    n8011[201] = 44'b00000000000000000000000000000000000000001001;
    n8011[200] = 44'b00000000000000000000000000000000000000000000;
    n8011[199] = 44'b00001011000000010000000100011101000110110001;
    n8011[198] = 44'b00000000000000000000000000000000000000000000;
    n8011[197] = 44'b00001010000000010000000100011100000110110001;
    n8011[196] = 44'b00001010000000010000000100011100000110110001;
    n8011[195] = 44'b00000000000000000000000000000000000000000000;
    n8011[194] = 44'b00000000000000000000000000000000000000000000;
    n8011[193] = 44'b00000000000000000000000000000000000000000000;
    n8011[192] = 44'b00000000000000000000000000000000000000000000;
    n8011[191] = 44'b00000000000000000000000000000000000000000000;
    n8011[190] = 44'b00000000000000000000000000000000000000000000;
    n8011[189] = 44'b00000000000000000000000000000000000000000000;
    n8011[188] = 44'b00000000000000000000000000000000000000000000;
    n8011[187] = 44'b00000000000000000000000000000000000000000000;
    n8011[186] = 44'b00000000000000000000000000000000000000000000;
    n8011[185] = 44'b00000000000000000000000000000000000000000000;
    n8011[184] = 44'b00000000000000000000000000000000000000000000;
    n8011[183] = 44'b00000000000000000000000000000000000000000000;
    n8011[182] = 44'b00000000000000000000000000000000000000000000;
    n8011[181] = 44'b00000000000000000000000000000000000000000000;
    n8011[180] = 44'b00000000000000000000000000000000000000000000;
    n8011[179] = 44'b00000000000000000000000000000000000000000000;
    n8011[178] = 44'b00000000000000000000000000000000000000000000;
    n8011[177] = 44'b00000000000000000000000000000000000000000000;
    n8011[176] = 44'b00000000000000000000010010000001010011101001;
    n8011[175] = 44'b00000000000000000000000000000000000000000000;
    n8011[174] = 44'b00000000000000000000000000000000000000000000;
    n8011[173] = 44'b00000000000000000000000000000000000000000000;
    n8011[172] = 44'b00000000000000000000000000000000000000000000;
    n8011[171] = 44'b00000000000000000000000000000000000000000000;
    n8011[170] = 44'b00000000000000100000000010000001010011111010;
    n8011[169] = 44'b00100000000000000000000000000000000000001001;
    n8011[168] = 44'b00000000001001100000001000000001010011111110;
    n8011[167] = 44'b00000000000000000000000000000000000000000000;
    n8011[166] = 44'b00000000000000000000000000000000000000000000;
    n8011[165] = 44'b00000000000000000000000000000000000000000000;
    n8011[164] = 44'b00000000000000000000000000000000000000000000;
    n8011[163] = 44'b00000000000000000000000000000000000000000000;
    n8011[162] = 44'b00000000000000000000000000000000000000000000;
    n8011[161] = 44'b00000000000000000000000000000000000000000000;
    n8011[160] = 44'b00000000000000000000000000000000000000000000;
    n8011[159] = 44'b00000000000000000000000000000000000000000000;
    n8011[158] = 44'b00000000000000000000000000000000000000000000;
    n8011[157] = 44'b00000000000000000000000000000000000000000000;
    n8011[156] = 44'b00000000000000000000000000000000000000000000;
    n8011[155] = 44'b00000000000000000000000000000000000000000000;
    n8011[154] = 44'b00000000000000000000000000000000000000000000;
    n8011[153] = 44'b00000000000000000000000000000000000000000000;
    n8011[152] = 44'b00000000000000000000000000000000000000000000;
    n8011[151] = 44'b00000000000000000000000000000000000000000000;
    n8011[150] = 44'b00000000000000000000000000000000000000000000;
    n8011[149] = 44'b00000000000000000000000000000000000000000000;
    n8011[148] = 44'b00000000000000000000000000000000000000000000;
    n8011[147] = 44'b00000000000000000000000000000000000000000000;
    n8011[146] = 44'b00000000000000000000000000000000000000000000;
    n8011[145] = 44'b00000000000000000000000000000000000000000000;
    n8011[144] = 44'b00000000000000000000010010000001010011101001;
    n8011[143] = 44'b00000000000000000000000000000000000000000000;
    n8011[142] = 44'b00000000000000000000000000000000000000000000;
    n8011[141] = 44'b00000000000000000000000000000000000000000000;
    n8011[140] = 44'b00000000000000000000000000000000000000000000;
    n8011[139] = 44'b00000000000000000000000000000000000000000000;
    n8011[138] = 44'b00000000000010000000000010000001010011111010;
    n8011[137] = 44'b00000000000000000000000000000000000000000000;
    n8011[136] = 44'b00000000000001100000001000000001010011111110;
    n8011[135] = 44'b00000000000000000000000000000000000000000000;
    n8011[134] = 44'b00000000000000000000000000000000000000000000;
    n8011[133] = 44'b00001000000000000000000100011100000011000001;
    n8011[132] = 44'b00001000000000000000000100011100000011000001;
    n8011[131] = 44'b00000000000000000000000000000000000000000000;
    n8011[130] = 44'b00000000000000000000000000000000000000000000;
    n8011[129] = 44'b00000000000000000000000000000000000000000000;
    n8011[128] = 44'b00000000000000000000000000000000000000000000;
    n8011[127] = 44'b00000000000000000000000000000000000000000000;
    n8011[126] = 44'b00000000000000000000000000000000000000000000;
    n8011[125] = 44'b00000000000000000000000000000000000000000000;
    n8011[124] = 44'b00000000000000000000000000000000000000000000;
    n8011[123] = 44'b00000000000000000000000000000000000000000000;
    n8011[122] = 44'b00000000000000000000000000000000000000000000;
    n8011[121] = 44'b00000000000000000000000000000000000000000000;
    n8011[120] = 44'b00000000000000000000000000000000000000000000;
    n8011[119] = 44'b00000000000000000000000000000000000000000000;
    n8011[118] = 44'b00001000000000000000000010000001001010110001;
    n8011[117] = 44'b00000000000000000000000000000000000000000000;
    n8011[116] = 44'b00001001000000000000000010000001001010110001;
    n8011[115] = 44'b00000000000000000000000000000000000000000000;
    n8011[114] = 44'b00000000000000000000000000000000000000000000;
    n8011[113] = 44'b00000000000000000000000000000000000000000000;
    n8011[112] = 44'b00000000000000000000010010000001010011101001;
    n8011[111] = 44'b00000000000000000000000000000000000000000000;
    n8011[110] = 44'b00000000000000000000000000000000000000000000;
    n8011[109] = 44'b00000000000000000000000000000000000000000000;
    n8011[108] = 44'b00000000000000000000000000000000000000000000;
    n8011[107] = 44'b00000000000000000000000000000000000000000000;
    n8011[106] = 44'b00000000000001100000000000010001010100000010;
    n8011[105] = 44'b00000000000101000000000000010001010100000010;
    n8011[104] = 44'b00000000000000000000000000000000000000000000;
    n8011[103] = 44'b00000000000000000000000000000000000000000000;
    n8011[102] = 44'b00000000000000000000000000000000000000000000;
    n8011[101] = 44'b00001000000001000000000100010000000010111001;
    n8011[100] = 44'b00000000000000000000000000000000000000000000;
    n8011[99] = 44'b00000000000000000000000000000000000000000000;
    n8011[98] = 44'b00000000000000000000000000000000000000000000;
    n8011[97] = 44'b00000000000000000000000000000000000000000000;
    n8011[96] = 44'b00000000000000000000000000000000000000000000;
    n8011[95] = 44'b00000000000000000000000000000000000000000000;
    n8011[94] = 44'b00000000000000000000000000000000000000000000;
    n8011[93] = 44'b00000000000000000000000000000000000000000000;
    n8011[92] = 44'b00000000000000000000000000000000000000000000;
    n8011[91] = 44'b00000000000000000000000000000000000000000000;
    n8011[90] = 44'b00000000000000000000000000000000000000000000;
    n8011[89] = 44'b00000000000000000000000000000000000000000000;
    n8011[88] = 44'b00000000000000000000000000000000000000000000;
    n8011[87] = 44'b00000000000000000000000000000000000000000000;
    n8011[86] = 44'b00001010000000000000000010000001001010110001;
    n8011[85] = 44'b00000000000000000000000000000000000000000000;
    n8011[84] = 44'b00001011000000000000000010000001001010110001;
    n8011[83] = 44'b00000000000000000000000000000000000000000000;
    n8011[82] = 44'b00000000000000000000000000000000000000000000;
    n8011[81] = 44'b00000000000000000000000000000000000000000000;
    n8011[80] = 44'b00000000000000000000010010000001010011101001;
    n8011[79] = 44'b00000000000000000000000000000000000000000000;
    n8011[78] = 44'b00000000000000000000000000000000000000000000;
    n8011[77] = 44'b00000000000000000000000000000000000000000000;
    n8011[76] = 44'b00000000000000000000000000000000000000000000;
    n8011[75] = 44'b00000000000000000000000000000000000000000000;
    n8011[74] = 44'b00000000000001000000000000010001010100000010;
    n8011[73] = 44'b00000000000000000000000000000000000000000000;
    n8011[72] = 44'b00000000000000000000000000000000000000000000;
    n8011[71] = 44'b00000000000000000000000000000000000000000000;
    n8011[70] = 44'b00000000000000000000000000000000000000000000;
    n8011[69] = 44'b00001000000000100000000100010000000010111001;
    n8011[68] = 44'b00000000000000000000000000000000000000000000;
    n8011[67] = 44'b00000000000000000000000000000000000000000000;
    n8011[66] = 44'b00000000000000000000000000000000000000000000;
    n8011[65] = 44'b00000000000000000000000000000000000000000000;
    n8011[64] = 44'b00000000000000000000000000000000000000000000;
    n8011[63] = 44'b00000000000000000000000000000000000000000000;
    n8011[62] = 44'b00000000000000000000000000000000000000000000;
    n8011[61] = 44'b00000000000000000000000000000000000000000000;
    n8011[60] = 44'b00000000000000000000000000000000000000000000;
    n8011[59] = 44'b00000000000000000000000000000000000000000000;
    n8011[58] = 44'b00000000000000000000000000000000000000000000;
    n8011[57] = 44'b00000000000000000000000000000000000000000000;
    n8011[56] = 44'b00000000000000000000000000000000000000000000;
    n8011[55] = 44'b00000000000000000000000000000000000000000000;
    n8011[54] = 44'b00001000000000000000000010000001001010101001;
    n8011[53] = 44'b00000000000000000000000000000000000000000000;
    n8011[52] = 44'b00001001000000000000000010000001001010101001;
    n8011[51] = 44'b00000000000000000000000000000000000000000000;
    n8011[50] = 44'b00000000000000000000000000000000000000000000;
    n8011[49] = 44'b00000000000000000000000000000000000000000000;
    n8011[48] = 44'b00000000000000000000010010000001010011101001;
    n8011[47] = 44'b00000000000000000000000000000000000000000000;
    n8011[46] = 44'b00000000000000000000000000000000000000000000;
    n8011[45] = 44'b00000000000000000000000000000000000000000000;
    n8011[44] = 44'b00000000000000000000000000000000000000000000;
    n8011[43] = 44'b00000000000000000000000000000000000000000000;
    n8011[42] = 44'b00000000000000100000000000010001010100000010;
    n8011[41] = 44'b00100000000000000000000000000000000011011001;
    n8011[40] = 44'b00000000000001100000000001000001010100000110;
    n8011[39] = 44'b00000000000000000000000000000000000000000000;
    n8011[38] = 44'b00000000000000000000000000000000000000000000;
    n8011[37] = 44'b00001000000001100000000100010000000010111001;
    n8011[36] = 44'b00000000000000000000000000000000000000000000;
    n8011[35] = 44'b00000000000000000000000000000000000000000000;
    n8011[34] = 44'b00000000000000000000000000000000000000000000;
    n8011[33] = 44'b00000000000000000000000000000000000000000000;
    n8011[32] = 44'b00000000000000000000000000000000000000000000;
    n8011[31] = 44'b00000000000000000000000000000000000000000000;
    n8011[30] = 44'b00000000000000000000000000000000000000000000;
    n8011[29] = 44'b00000000000000000000000000000000000000000000;
    n8011[28] = 44'b00000000000000000000000000000000000000000000;
    n8011[27] = 44'b00000000000000000000000000000000000000000000;
    n8011[26] = 44'b00000000000000000000000000000000000000000000;
    n8011[25] = 44'b00000000000000000000000000000000000000000000;
    n8011[24] = 44'b00000000000000000000000000000000000000000000;
    n8011[23] = 44'b00000000000000000000000000000000000000000000;
    n8011[22] = 44'b00001010000000000000000010000001001010101001;
    n8011[21] = 44'b00000000000000000000000000000000000000000000;
    n8011[20] = 44'b00001011000000000000000010000001001010101001;
    n8011[19] = 44'b00000000000000000000000000000000000000000000;
    n8011[18] = 44'b00000000000000000000000000000000000000000000;
    n8011[17] = 44'b00000000000000000000000000000000000000000000;
    n8011[16] = 44'b00000000000000000000010010000001010011101001;
    n8011[15] = 44'b00000000000000000000000000000000000000000000;
    n8011[14] = 44'b00000000000000000000000000000000000000000000;
    n8011[13] = 44'b00000000000000000000000000000000000000000000;
    n8011[12] = 44'b00000000000000000000000000000000000000000000;
    n8011[11] = 44'b00000000000000000000000000000000000000000000;
    n8011[10] = 44'b00000000000010000000000000010001010100000010;
    n8011[9] = 44'b00000000000000000000000000000001010010100010;
    n8011[8] = 44'b00000000000000000000000000000000000000000000;
    n8011[7] = 44'b00000000000000000000000000000000000000000000;
    n8011[6] = 44'b00000000000000000000000000000000000000000000;
    n8011[5] = 44'b00000000000000000000000000000000000000000000;
    n8011[4] = 44'b00000000000000000000000000000000000000000000;
    n8011[3] = 44'b00000000000000000000000000000000000000000000;
    n8011[2] = 44'b00000000000000000000000000000000000000000000;
    n8011[1] = 44'b00000000000000000000000000000000000000000000;
    n8011[0] = 44'b00000000000000000000000000000000000000000000;
    end
  assign n8012_data = n8011[n7465_o];
  /* decode1.vhdl:598:44  */
  /* decode1.vhdl:598:43  */
  reg n8013[1023:0] ; // memory
  initial begin
    n8013[1023] = 1'b1;
    n8013[1022] = 1'b0;
    n8013[1021] = 1'b0;
    n8013[1020] = 1'b0;
    n8013[1019] = 1'b0;
    n8013[1018] = 1'b0;
    n8013[1017] = 1'b0;
    n8013[1016] = 1'b0;
    n8013[1015] = 1'b0;
    n8013[1014] = 1'b0;
    n8013[1013] = 1'b0;
    n8013[1012] = 1'b0;
    n8013[1011] = 1'b0;
    n8013[1010] = 1'b0;
    n8013[1009] = 1'b0;
    n8013[1008] = 1'b0;
    n8013[1007] = 1'b0;
    n8013[1006] = 1'b0;
    n8013[1005] = 1'b0;
    n8013[1004] = 1'b0;
    n8013[1003] = 1'b0;
    n8013[1002] = 1'b0;
    n8013[1001] = 1'b0;
    n8013[1000] = 1'b0;
    n8013[999] = 1'b0;
    n8013[998] = 1'b0;
    n8013[997] = 1'b0;
    n8013[996] = 1'b0;
    n8013[995] = 1'b0;
    n8013[994] = 1'b0;
    n8013[993] = 1'b0;
    n8013[992] = 1'b0;
    n8013[991] = 1'b0;
    n8013[990] = 1'b1;
    n8013[989] = 1'b0;
    n8013[988] = 1'b0;
    n8013[987] = 1'b1;
    n8013[986] = 1'b0;
    n8013[985] = 1'b1;
    n8013[984] = 1'b1;
    n8013[983] = 1'b1;
    n8013[982] = 1'b1;
    n8013[981] = 1'b0;
    n8013[980] = 1'b0;
    n8013[979] = 1'b0;
    n8013[978] = 1'b1;
    n8013[977] = 1'b1;
    n8013[976] = 1'b0;
    n8013[975] = 1'b0;
    n8013[974] = 1'b0;
    n8013[973] = 1'b0;
    n8013[972] = 1'b0;
    n8013[971] = 1'b0;
    n8013[970] = 1'b0;
    n8013[969] = 1'b0;
    n8013[968] = 1'b0;
    n8013[967] = 1'b0;
    n8013[966] = 1'b0;
    n8013[965] = 1'b0;
    n8013[964] = 1'b0;
    n8013[963] = 1'b0;
    n8013[962] = 1'b0;
    n8013[961] = 1'b0;
    n8013[960] = 1'b0;
    n8013[959] = 1'b1;
    n8013[958] = 1'b1;
    n8013[957] = 1'b1;
    n8013[956] = 1'b1;
    n8013[955] = 1'b1;
    n8013[954] = 1'b1;
    n8013[953] = 1'b1;
    n8013[952] = 1'b1;
    n8013[951] = 1'b1;
    n8013[950] = 1'b1;
    n8013[949] = 1'b1;
    n8013[948] = 1'b1;
    n8013[947] = 1'b1;
    n8013[946] = 1'b1;
    n8013[945] = 1'b1;
    n8013[944] = 1'b1;
    n8013[943] = 1'b1;
    n8013[942] = 1'b1;
    n8013[941] = 1'b1;
    n8013[940] = 1'b1;
    n8013[939] = 1'b1;
    n8013[938] = 1'b1;
    n8013[937] = 1'b1;
    n8013[936] = 1'b1;
    n8013[935] = 1'b1;
    n8013[934] = 1'b1;
    n8013[933] = 1'b1;
    n8013[932] = 1'b1;
    n8013[931] = 1'b1;
    n8013[930] = 1'b1;
    n8013[929] = 1'b1;
    n8013[928] = 1'b1;
    n8013[927] = 1'b0;
    n8013[926] = 1'b0;
    n8013[925] = 1'b0;
    n8013[924] = 1'b0;
    n8013[923] = 1'b0;
    n8013[922] = 1'b0;
    n8013[921] = 1'b0;
    n8013[920] = 1'b0;
    n8013[919] = 1'b0;
    n8013[918] = 1'b0;
    n8013[917] = 1'b0;
    n8013[916] = 1'b0;
    n8013[915] = 1'b0;
    n8013[914] = 1'b0;
    n8013[913] = 1'b0;
    n8013[912] = 1'b0;
    n8013[911] = 1'b0;
    n8013[910] = 1'b0;
    n8013[909] = 1'b0;
    n8013[908] = 1'b0;
    n8013[907] = 1'b0;
    n8013[906] = 1'b0;
    n8013[905] = 1'b0;
    n8013[904] = 1'b0;
    n8013[903] = 1'b0;
    n8013[902] = 1'b0;
    n8013[901] = 1'b0;
    n8013[900] = 1'b0;
    n8013[899] = 1'b0;
    n8013[898] = 1'b0;
    n8013[897] = 1'b0;
    n8013[896] = 1'b0;
    n8013[895] = 1'b0;
    n8013[894] = 1'b0;
    n8013[893] = 1'b0;
    n8013[892] = 1'b0;
    n8013[891] = 1'b0;
    n8013[890] = 1'b0;
    n8013[889] = 1'b0;
    n8013[888] = 1'b0;
    n8013[887] = 1'b0;
    n8013[886] = 1'b0;
    n8013[885] = 1'b0;
    n8013[884] = 1'b0;
    n8013[883] = 1'b0;
    n8013[882] = 1'b0;
    n8013[881] = 1'b0;
    n8013[880] = 1'b0;
    n8013[879] = 1'b0;
    n8013[878] = 1'b0;
    n8013[877] = 1'b0;
    n8013[876] = 1'b0;
    n8013[875] = 1'b0;
    n8013[874] = 1'b0;
    n8013[873] = 1'b0;
    n8013[872] = 1'b0;
    n8013[871] = 1'b0;
    n8013[870] = 1'b0;
    n8013[869] = 1'b0;
    n8013[868] = 1'b0;
    n8013[867] = 1'b0;
    n8013[866] = 1'b0;
    n8013[865] = 1'b0;
    n8013[864] = 1'b0;
    n8013[863] = 1'b0;
    n8013[862] = 1'b0;
    n8013[861] = 1'b0;
    n8013[860] = 1'b0;
    n8013[859] = 1'b0;
    n8013[858] = 1'b0;
    n8013[857] = 1'b0;
    n8013[856] = 1'b0;
    n8013[855] = 1'b0;
    n8013[854] = 1'b0;
    n8013[853] = 1'b0;
    n8013[852] = 1'b0;
    n8013[851] = 1'b0;
    n8013[850] = 1'b0;
    n8013[849] = 1'b0;
    n8013[848] = 1'b0;
    n8013[847] = 1'b0;
    n8013[846] = 1'b0;
    n8013[845] = 1'b0;
    n8013[844] = 1'b0;
    n8013[843] = 1'b0;
    n8013[842] = 1'b0;
    n8013[841] = 1'b0;
    n8013[840] = 1'b0;
    n8013[839] = 1'b0;
    n8013[838] = 1'b0;
    n8013[837] = 1'b0;
    n8013[836] = 1'b0;
    n8013[835] = 1'b0;
    n8013[834] = 1'b0;
    n8013[833] = 1'b0;
    n8013[832] = 1'b0;
    n8013[831] = 1'b0;
    n8013[830] = 1'b0;
    n8013[829] = 1'b0;
    n8013[828] = 1'b0;
    n8013[827] = 1'b0;
    n8013[826] = 1'b0;
    n8013[825] = 1'b0;
    n8013[824] = 1'b0;
    n8013[823] = 1'b0;
    n8013[822] = 1'b0;
    n8013[821] = 1'b0;
    n8013[820] = 1'b0;
    n8013[819] = 1'b0;
    n8013[818] = 1'b0;
    n8013[817] = 1'b0;
    n8013[816] = 1'b0;
    n8013[815] = 1'b0;
    n8013[814] = 1'b0;
    n8013[813] = 1'b0;
    n8013[812] = 1'b0;
    n8013[811] = 1'b0;
    n8013[810] = 1'b0;
    n8013[809] = 1'b0;
    n8013[808] = 1'b0;
    n8013[807] = 1'b0;
    n8013[806] = 1'b0;
    n8013[805] = 1'b0;
    n8013[804] = 1'b0;
    n8013[803] = 1'b0;
    n8013[802] = 1'b0;
    n8013[801] = 1'b0;
    n8013[800] = 1'b0;
    n8013[799] = 1'b0;
    n8013[798] = 1'b0;
    n8013[797] = 1'b0;
    n8013[796] = 1'b0;
    n8013[795] = 1'b0;
    n8013[794] = 1'b0;
    n8013[793] = 1'b0;
    n8013[792] = 1'b0;
    n8013[791] = 1'b0;
    n8013[790] = 1'b0;
    n8013[789] = 1'b0;
    n8013[788] = 1'b0;
    n8013[787] = 1'b0;
    n8013[786] = 1'b0;
    n8013[785] = 1'b0;
    n8013[784] = 1'b0;
    n8013[783] = 1'b0;
    n8013[782] = 1'b0;
    n8013[781] = 1'b0;
    n8013[780] = 1'b0;
    n8013[779] = 1'b0;
    n8013[778] = 1'b0;
    n8013[777] = 1'b0;
    n8013[776] = 1'b0;
    n8013[775] = 1'b0;
    n8013[774] = 1'b0;
    n8013[773] = 1'b0;
    n8013[772] = 1'b0;
    n8013[771] = 1'b0;
    n8013[770] = 1'b0;
    n8013[769] = 1'b0;
    n8013[768] = 1'b0;
    n8013[767] = 1'b0;
    n8013[766] = 1'b0;
    n8013[765] = 1'b0;
    n8013[764] = 1'b0;
    n8013[763] = 1'b0;
    n8013[762] = 1'b0;
    n8013[761] = 1'b0;
    n8013[760] = 1'b0;
    n8013[759] = 1'b0;
    n8013[758] = 1'b0;
    n8013[757] = 1'b0;
    n8013[756] = 1'b0;
    n8013[755] = 1'b0;
    n8013[754] = 1'b0;
    n8013[753] = 1'b0;
    n8013[752] = 1'b0;
    n8013[751] = 1'b0;
    n8013[750] = 1'b0;
    n8013[749] = 1'b0;
    n8013[748] = 1'b0;
    n8013[747] = 1'b0;
    n8013[746] = 1'b0;
    n8013[745] = 1'b0;
    n8013[744] = 1'b0;
    n8013[743] = 1'b0;
    n8013[742] = 1'b0;
    n8013[741] = 1'b0;
    n8013[740] = 1'b0;
    n8013[739] = 1'b0;
    n8013[738] = 1'b0;
    n8013[737] = 1'b0;
    n8013[736] = 1'b0;
    n8013[735] = 1'b0;
    n8013[734] = 1'b0;
    n8013[733] = 1'b0;
    n8013[732] = 1'b0;
    n8013[731] = 1'b0;
    n8013[730] = 1'b0;
    n8013[729] = 1'b0;
    n8013[728] = 1'b0;
    n8013[727] = 1'b0;
    n8013[726] = 1'b0;
    n8013[725] = 1'b0;
    n8013[724] = 1'b0;
    n8013[723] = 1'b0;
    n8013[722] = 1'b0;
    n8013[721] = 1'b0;
    n8013[720] = 1'b0;
    n8013[719] = 1'b0;
    n8013[718] = 1'b0;
    n8013[717] = 1'b0;
    n8013[716] = 1'b0;
    n8013[715] = 1'b0;
    n8013[714] = 1'b0;
    n8013[713] = 1'b0;
    n8013[712] = 1'b0;
    n8013[711] = 1'b0;
    n8013[710] = 1'b0;
    n8013[709] = 1'b0;
    n8013[708] = 1'b0;
    n8013[707] = 1'b0;
    n8013[706] = 1'b0;
    n8013[705] = 1'b0;
    n8013[704] = 1'b0;
    n8013[703] = 1'b0;
    n8013[702] = 1'b0;
    n8013[701] = 1'b0;
    n8013[700] = 1'b0;
    n8013[699] = 1'b0;
    n8013[698] = 1'b0;
    n8013[697] = 1'b0;
    n8013[696] = 1'b0;
    n8013[695] = 1'b0;
    n8013[694] = 1'b0;
    n8013[693] = 1'b0;
    n8013[692] = 1'b0;
    n8013[691] = 1'b0;
    n8013[690] = 1'b0;
    n8013[689] = 1'b0;
    n8013[688] = 1'b0;
    n8013[687] = 1'b0;
    n8013[686] = 1'b0;
    n8013[685] = 1'b0;
    n8013[684] = 1'b0;
    n8013[683] = 1'b0;
    n8013[682] = 1'b0;
    n8013[681] = 1'b0;
    n8013[680] = 1'b0;
    n8013[679] = 1'b0;
    n8013[678] = 1'b0;
    n8013[677] = 1'b0;
    n8013[676] = 1'b0;
    n8013[675] = 1'b0;
    n8013[674] = 1'b0;
    n8013[673] = 1'b0;
    n8013[672] = 1'b0;
    n8013[671] = 1'b0;
    n8013[670] = 1'b0;
    n8013[669] = 1'b0;
    n8013[668] = 1'b0;
    n8013[667] = 1'b0;
    n8013[666] = 1'b0;
    n8013[665] = 1'b0;
    n8013[664] = 1'b0;
    n8013[663] = 1'b0;
    n8013[662] = 1'b0;
    n8013[661] = 1'b0;
    n8013[660] = 1'b0;
    n8013[659] = 1'b0;
    n8013[658] = 1'b0;
    n8013[657] = 1'b0;
    n8013[656] = 1'b0;
    n8013[655] = 1'b0;
    n8013[654] = 1'b0;
    n8013[653] = 1'b0;
    n8013[652] = 1'b0;
    n8013[651] = 1'b0;
    n8013[650] = 1'b0;
    n8013[649] = 1'b0;
    n8013[648] = 1'b0;
    n8013[647] = 1'b0;
    n8013[646] = 1'b0;
    n8013[645] = 1'b0;
    n8013[644] = 1'b0;
    n8013[643] = 1'b0;
    n8013[642] = 1'b0;
    n8013[641] = 1'b0;
    n8013[640] = 1'b0;
    n8013[639] = 1'b0;
    n8013[638] = 1'b0;
    n8013[637] = 1'b0;
    n8013[636] = 1'b0;
    n8013[635] = 1'b0;
    n8013[634] = 1'b0;
    n8013[633] = 1'b0;
    n8013[632] = 1'b0;
    n8013[631] = 1'b0;
    n8013[630] = 1'b0;
    n8013[629] = 1'b0;
    n8013[628] = 1'b0;
    n8013[627] = 1'b0;
    n8013[626] = 1'b0;
    n8013[625] = 1'b0;
    n8013[624] = 1'b0;
    n8013[623] = 1'b0;
    n8013[622] = 1'b0;
    n8013[621] = 1'b0;
    n8013[620] = 1'b0;
    n8013[619] = 1'b0;
    n8013[618] = 1'b0;
    n8013[617] = 1'b0;
    n8013[616] = 1'b0;
    n8013[615] = 1'b0;
    n8013[614] = 1'b0;
    n8013[613] = 1'b0;
    n8013[612] = 1'b0;
    n8013[611] = 1'b0;
    n8013[610] = 1'b0;
    n8013[609] = 1'b0;
    n8013[608] = 1'b0;
    n8013[607] = 1'b0;
    n8013[606] = 1'b0;
    n8013[605] = 1'b0;
    n8013[604] = 1'b0;
    n8013[603] = 1'b0;
    n8013[602] = 1'b0;
    n8013[601] = 1'b0;
    n8013[600] = 1'b0;
    n8013[599] = 1'b0;
    n8013[598] = 1'b0;
    n8013[597] = 1'b0;
    n8013[596] = 1'b0;
    n8013[595] = 1'b0;
    n8013[594] = 1'b0;
    n8013[593] = 1'b0;
    n8013[592] = 1'b0;
    n8013[591] = 1'b0;
    n8013[590] = 1'b0;
    n8013[589] = 1'b0;
    n8013[588] = 1'b0;
    n8013[587] = 1'b0;
    n8013[586] = 1'b0;
    n8013[585] = 1'b0;
    n8013[584] = 1'b0;
    n8013[583] = 1'b0;
    n8013[582] = 1'b0;
    n8013[581] = 1'b0;
    n8013[580] = 1'b0;
    n8013[579] = 1'b0;
    n8013[578] = 1'b0;
    n8013[577] = 1'b0;
    n8013[576] = 1'b0;
    n8013[575] = 1'b0;
    n8013[574] = 1'b0;
    n8013[573] = 1'b0;
    n8013[572] = 1'b0;
    n8013[571] = 1'b0;
    n8013[570] = 1'b0;
    n8013[569] = 1'b0;
    n8013[568] = 1'b0;
    n8013[567] = 1'b0;
    n8013[566] = 1'b0;
    n8013[565] = 1'b0;
    n8013[564] = 1'b0;
    n8013[563] = 1'b0;
    n8013[562] = 1'b0;
    n8013[561] = 1'b0;
    n8013[560] = 1'b0;
    n8013[559] = 1'b0;
    n8013[558] = 1'b0;
    n8013[557] = 1'b0;
    n8013[556] = 1'b0;
    n8013[555] = 1'b0;
    n8013[554] = 1'b0;
    n8013[553] = 1'b0;
    n8013[552] = 1'b0;
    n8013[551] = 1'b0;
    n8013[550] = 1'b0;
    n8013[549] = 1'b0;
    n8013[548] = 1'b0;
    n8013[547] = 1'b0;
    n8013[546] = 1'b0;
    n8013[545] = 1'b0;
    n8013[544] = 1'b0;
    n8013[543] = 1'b0;
    n8013[542] = 1'b0;
    n8013[541] = 1'b0;
    n8013[540] = 1'b0;
    n8013[539] = 1'b0;
    n8013[538] = 1'b0;
    n8013[537] = 1'b0;
    n8013[536] = 1'b0;
    n8013[535] = 1'b0;
    n8013[534] = 1'b0;
    n8013[533] = 1'b0;
    n8013[532] = 1'b0;
    n8013[531] = 1'b0;
    n8013[530] = 1'b0;
    n8013[529] = 1'b0;
    n8013[528] = 1'b0;
    n8013[527] = 1'b0;
    n8013[526] = 1'b0;
    n8013[525] = 1'b0;
    n8013[524] = 1'b0;
    n8013[523] = 1'b0;
    n8013[522] = 1'b0;
    n8013[521] = 1'b0;
    n8013[520] = 1'b0;
    n8013[519] = 1'b0;
    n8013[518] = 1'b0;
    n8013[517] = 1'b0;
    n8013[516] = 1'b0;
    n8013[515] = 1'b0;
    n8013[514] = 1'b0;
    n8013[513] = 1'b0;
    n8013[512] = 1'b0;
    n8013[511] = 1'b1;
    n8013[510] = 1'b0;
    n8013[509] = 1'b0;
    n8013[508] = 1'b0;
    n8013[507] = 1'b0;
    n8013[506] = 1'b0;
    n8013[505] = 1'b0;
    n8013[504] = 1'b0;
    n8013[503] = 1'b0;
    n8013[502] = 1'b0;
    n8013[501] = 1'b0;
    n8013[500] = 1'b0;
    n8013[499] = 1'b0;
    n8013[498] = 1'b0;
    n8013[497] = 1'b0;
    n8013[496] = 1'b0;
    n8013[495] = 1'b1;
    n8013[494] = 1'b1;
    n8013[493] = 1'b0;
    n8013[492] = 1'b0;
    n8013[491] = 1'b0;
    n8013[490] = 1'b0;
    n8013[489] = 1'b0;
    n8013[488] = 1'b0;
    n8013[487] = 1'b0;
    n8013[486] = 1'b0;
    n8013[485] = 1'b0;
    n8013[484] = 1'b0;
    n8013[483] = 1'b0;
    n8013[482] = 1'b0;
    n8013[481] = 1'b0;
    n8013[480] = 1'b0;
    n8013[479] = 1'b0;
    n8013[478] = 1'b0;
    n8013[477] = 1'b0;
    n8013[476] = 1'b0;
    n8013[475] = 1'b0;
    n8013[474] = 1'b0;
    n8013[473] = 1'b0;
    n8013[472] = 1'b0;
    n8013[471] = 1'b0;
    n8013[470] = 1'b0;
    n8013[469] = 1'b0;
    n8013[468] = 1'b0;
    n8013[467] = 1'b0;
    n8013[466] = 1'b0;
    n8013[465] = 1'b0;
    n8013[464] = 1'b0;
    n8013[463] = 1'b0;
    n8013[462] = 1'b0;
    n8013[461] = 1'b0;
    n8013[460] = 1'b0;
    n8013[459] = 1'b0;
    n8013[458] = 1'b0;
    n8013[457] = 1'b0;
    n8013[456] = 1'b0;
    n8013[455] = 1'b0;
    n8013[454] = 1'b0;
    n8013[453] = 1'b0;
    n8013[452] = 1'b0;
    n8013[451] = 1'b0;
    n8013[450] = 1'b0;
    n8013[449] = 1'b0;
    n8013[448] = 1'b0;
    n8013[447] = 1'b1;
    n8013[446] = 1'b0;
    n8013[445] = 1'b0;
    n8013[444] = 1'b0;
    n8013[443] = 1'b0;
    n8013[442] = 1'b0;
    n8013[441] = 1'b0;
    n8013[440] = 1'b0;
    n8013[439] = 1'b0;
    n8013[438] = 1'b0;
    n8013[437] = 1'b0;
    n8013[436] = 1'b0;
    n8013[435] = 1'b0;
    n8013[434] = 1'b0;
    n8013[433] = 1'b0;
    n8013[432] = 1'b0;
    n8013[431] = 1'b0;
    n8013[430] = 1'b0;
    n8013[429] = 1'b0;
    n8013[428] = 1'b0;
    n8013[427] = 1'b0;
    n8013[426] = 1'b0;
    n8013[425] = 1'b0;
    n8013[424] = 1'b0;
    n8013[423] = 1'b0;
    n8013[422] = 1'b0;
    n8013[421] = 1'b0;
    n8013[420] = 1'b0;
    n8013[419] = 1'b0;
    n8013[418] = 1'b0;
    n8013[417] = 1'b0;
    n8013[416] = 1'b0;
    n8013[415] = 1'b0;
    n8013[414] = 1'b0;
    n8013[413] = 1'b0;
    n8013[412] = 1'b0;
    n8013[411] = 1'b0;
    n8013[410] = 1'b0;
    n8013[409] = 1'b0;
    n8013[408] = 1'b0;
    n8013[407] = 1'b0;
    n8013[406] = 1'b0;
    n8013[405] = 1'b0;
    n8013[404] = 1'b0;
    n8013[403] = 1'b0;
    n8013[402] = 1'b0;
    n8013[401] = 1'b0;
    n8013[400] = 1'b0;
    n8013[399] = 1'b0;
    n8013[398] = 1'b0;
    n8013[397] = 1'b0;
    n8013[396] = 1'b0;
    n8013[395] = 1'b0;
    n8013[394] = 1'b0;
    n8013[393] = 1'b0;
    n8013[392] = 1'b0;
    n8013[391] = 1'b0;
    n8013[390] = 1'b0;
    n8013[389] = 1'b0;
    n8013[388] = 1'b0;
    n8013[387] = 1'b0;
    n8013[386] = 1'b0;
    n8013[385] = 1'b0;
    n8013[384] = 1'b0;
    n8013[383] = 1'b0;
    n8013[382] = 1'b0;
    n8013[381] = 1'b0;
    n8013[380] = 1'b0;
    n8013[379] = 1'b0;
    n8013[378] = 1'b0;
    n8013[377] = 1'b0;
    n8013[376] = 1'b0;
    n8013[375] = 1'b0;
    n8013[374] = 1'b0;
    n8013[373] = 1'b0;
    n8013[372] = 1'b0;
    n8013[371] = 1'b0;
    n8013[370] = 1'b0;
    n8013[369] = 1'b0;
    n8013[368] = 1'b0;
    n8013[367] = 1'b0;
    n8013[366] = 1'b0;
    n8013[365] = 1'b0;
    n8013[364] = 1'b0;
    n8013[363] = 1'b0;
    n8013[362] = 1'b0;
    n8013[361] = 1'b0;
    n8013[360] = 1'b0;
    n8013[359] = 1'b0;
    n8013[358] = 1'b0;
    n8013[357] = 1'b0;
    n8013[356] = 1'b0;
    n8013[355] = 1'b0;
    n8013[354] = 1'b0;
    n8013[353] = 1'b0;
    n8013[352] = 1'b0;
    n8013[351] = 1'b0;
    n8013[350] = 1'b0;
    n8013[349] = 1'b0;
    n8013[348] = 1'b0;
    n8013[347] = 1'b0;
    n8013[346] = 1'b0;
    n8013[345] = 1'b0;
    n8013[344] = 1'b0;
    n8013[343] = 1'b0;
    n8013[342] = 1'b0;
    n8013[341] = 1'b0;
    n8013[340] = 1'b0;
    n8013[339] = 1'b0;
    n8013[338] = 1'b0;
    n8013[337] = 1'b0;
    n8013[336] = 1'b0;
    n8013[335] = 1'b0;
    n8013[334] = 1'b0;
    n8013[333] = 1'b0;
    n8013[332] = 1'b0;
    n8013[331] = 1'b0;
    n8013[330] = 1'b0;
    n8013[329] = 1'b0;
    n8013[328] = 1'b0;
    n8013[327] = 1'b0;
    n8013[326] = 1'b0;
    n8013[325] = 1'b0;
    n8013[324] = 1'b0;
    n8013[323] = 1'b0;
    n8013[322] = 1'b0;
    n8013[321] = 1'b0;
    n8013[320] = 1'b0;
    n8013[319] = 1'b0;
    n8013[318] = 1'b0;
    n8013[317] = 1'b0;
    n8013[316] = 1'b0;
    n8013[315] = 1'b1;
    n8013[314] = 1'b0;
    n8013[313] = 1'b0;
    n8013[312] = 1'b0;
    n8013[311] = 1'b0;
    n8013[310] = 1'b0;
    n8013[309] = 1'b0;
    n8013[308] = 1'b0;
    n8013[307] = 1'b0;
    n8013[306] = 1'b0;
    n8013[305] = 1'b0;
    n8013[304] = 1'b0;
    n8013[303] = 1'b0;
    n8013[302] = 1'b0;
    n8013[301] = 1'b0;
    n8013[300] = 1'b0;
    n8013[299] = 1'b0;
    n8013[298] = 1'b0;
    n8013[297] = 1'b0;
    n8013[296] = 1'b0;
    n8013[295] = 1'b0;
    n8013[294] = 1'b0;
    n8013[293] = 1'b0;
    n8013[292] = 1'b0;
    n8013[291] = 1'b0;
    n8013[290] = 1'b0;
    n8013[289] = 1'b0;
    n8013[288] = 1'b0;
    n8013[287] = 1'b0;
    n8013[286] = 1'b0;
    n8013[285] = 1'b0;
    n8013[284] = 1'b0;
    n8013[283] = 1'b0;
    n8013[282] = 1'b0;
    n8013[281] = 1'b0;
    n8013[280] = 1'b0;
    n8013[279] = 1'b0;
    n8013[278] = 1'b0;
    n8013[277] = 1'b0;
    n8013[276] = 1'b0;
    n8013[275] = 1'b0;
    n8013[274] = 1'b0;
    n8013[273] = 1'b0;
    n8013[272] = 1'b0;
    n8013[271] = 1'b0;
    n8013[270] = 1'b0;
    n8013[269] = 1'b0;
    n8013[268] = 1'b0;
    n8013[267] = 1'b0;
    n8013[266] = 1'b0;
    n8013[265] = 1'b0;
    n8013[264] = 1'b0;
    n8013[263] = 1'b0;
    n8013[262] = 1'b0;
    n8013[261] = 1'b0;
    n8013[260] = 1'b0;
    n8013[259] = 1'b0;
    n8013[258] = 1'b0;
    n8013[257] = 1'b0;
    n8013[256] = 1'b0;
    n8013[255] = 1'b0;
    n8013[254] = 1'b0;
    n8013[253] = 1'b0;
    n8013[252] = 1'b0;
    n8013[251] = 1'b0;
    n8013[250] = 1'b0;
    n8013[249] = 1'b0;
    n8013[248] = 1'b0;
    n8013[247] = 1'b0;
    n8013[246] = 1'b0;
    n8013[245] = 1'b0;
    n8013[244] = 1'b0;
    n8013[243] = 1'b0;
    n8013[242] = 1'b0;
    n8013[241] = 1'b0;
    n8013[240] = 1'b0;
    n8013[239] = 1'b0;
    n8013[238] = 1'b0;
    n8013[237] = 1'b0;
    n8013[236] = 1'b0;
    n8013[235] = 1'b0;
    n8013[234] = 1'b0;
    n8013[233] = 1'b0;
    n8013[232] = 1'b0;
    n8013[231] = 1'b0;
    n8013[230] = 1'b0;
    n8013[229] = 1'b0;
    n8013[228] = 1'b0;
    n8013[227] = 1'b0;
    n8013[226] = 1'b0;
    n8013[225] = 1'b0;
    n8013[224] = 1'b0;
    n8013[223] = 1'b0;
    n8013[222] = 1'b0;
    n8013[221] = 1'b0;
    n8013[220] = 1'b0;
    n8013[219] = 1'b0;
    n8013[218] = 1'b0;
    n8013[217] = 1'b0;
    n8013[216] = 1'b0;
    n8013[215] = 1'b0;
    n8013[214] = 1'b0;
    n8013[213] = 1'b0;
    n8013[212] = 1'b0;
    n8013[211] = 1'b0;
    n8013[210] = 1'b0;
    n8013[209] = 1'b0;
    n8013[208] = 1'b0;
    n8013[207] = 1'b0;
    n8013[206] = 1'b0;
    n8013[205] = 1'b0;
    n8013[204] = 1'b0;
    n8013[203] = 1'b0;
    n8013[202] = 1'b0;
    n8013[201] = 1'b0;
    n8013[200] = 1'b0;
    n8013[199] = 1'b0;
    n8013[198] = 1'b0;
    n8013[197] = 1'b0;
    n8013[196] = 1'b0;
    n8013[195] = 1'b0;
    n8013[194] = 1'b0;
    n8013[193] = 1'b0;
    n8013[192] = 1'b0;
    n8013[191] = 1'b0;
    n8013[190] = 1'b0;
    n8013[189] = 1'b0;
    n8013[188] = 1'b0;
    n8013[187] = 1'b0;
    n8013[186] = 1'b0;
    n8013[185] = 1'b0;
    n8013[184] = 1'b0;
    n8013[183] = 1'b0;
    n8013[182] = 1'b0;
    n8013[181] = 1'b0;
    n8013[180] = 1'b0;
    n8013[179] = 1'b0;
    n8013[178] = 1'b0;
    n8013[177] = 1'b0;
    n8013[176] = 1'b0;
    n8013[175] = 1'b0;
    n8013[174] = 1'b0;
    n8013[173] = 1'b0;
    n8013[172] = 1'b0;
    n8013[171] = 1'b0;
    n8013[170] = 1'b0;
    n8013[169] = 1'b0;
    n8013[168] = 1'b0;
    n8013[167] = 1'b0;
    n8013[166] = 1'b0;
    n8013[165] = 1'b0;
    n8013[164] = 1'b0;
    n8013[163] = 1'b0;
    n8013[162] = 1'b0;
    n8013[161] = 1'b0;
    n8013[160] = 1'b0;
    n8013[159] = 1'b0;
    n8013[158] = 1'b0;
    n8013[157] = 1'b0;
    n8013[156] = 1'b0;
    n8013[155] = 1'b0;
    n8013[154] = 1'b0;
    n8013[153] = 1'b0;
    n8013[152] = 1'b0;
    n8013[151] = 1'b0;
    n8013[150] = 1'b0;
    n8013[149] = 1'b0;
    n8013[148] = 1'b0;
    n8013[147] = 1'b0;
    n8013[146] = 1'b0;
    n8013[145] = 1'b0;
    n8013[144] = 1'b0;
    n8013[143] = 1'b0;
    n8013[142] = 1'b0;
    n8013[141] = 1'b0;
    n8013[140] = 1'b0;
    n8013[139] = 1'b0;
    n8013[138] = 1'b0;
    n8013[137] = 1'b0;
    n8013[136] = 1'b0;
    n8013[135] = 1'b0;
    n8013[134] = 1'b0;
    n8013[133] = 1'b0;
    n8013[132] = 1'b0;
    n8013[131] = 1'b0;
    n8013[130] = 1'b0;
    n8013[129] = 1'b0;
    n8013[128] = 1'b0;
    n8013[127] = 1'b0;
    n8013[126] = 1'b0;
    n8013[125] = 1'b0;
    n8013[124] = 1'b0;
    n8013[123] = 1'b0;
    n8013[122] = 1'b0;
    n8013[121] = 1'b0;
    n8013[120] = 1'b0;
    n8013[119] = 1'b0;
    n8013[118] = 1'b0;
    n8013[117] = 1'b0;
    n8013[116] = 1'b0;
    n8013[115] = 1'b0;
    n8013[114] = 1'b0;
    n8013[113] = 1'b0;
    n8013[112] = 1'b0;
    n8013[111] = 1'b0;
    n8013[110] = 1'b0;
    n8013[109] = 1'b0;
    n8013[108] = 1'b0;
    n8013[107] = 1'b0;
    n8013[106] = 1'b0;
    n8013[105] = 1'b0;
    n8013[104] = 1'b0;
    n8013[103] = 1'b0;
    n8013[102] = 1'b0;
    n8013[101] = 1'b0;
    n8013[100] = 1'b0;
    n8013[99] = 1'b0;
    n8013[98] = 1'b0;
    n8013[97] = 1'b0;
    n8013[96] = 1'b0;
    n8013[95] = 1'b0;
    n8013[94] = 1'b0;
    n8013[93] = 1'b0;
    n8013[92] = 1'b0;
    n8013[91] = 1'b0;
    n8013[90] = 1'b0;
    n8013[89] = 1'b0;
    n8013[88] = 1'b0;
    n8013[87] = 1'b0;
    n8013[86] = 1'b0;
    n8013[85] = 1'b0;
    n8013[84] = 1'b0;
    n8013[83] = 1'b0;
    n8013[82] = 1'b0;
    n8013[81] = 1'b0;
    n8013[80] = 1'b0;
    n8013[79] = 1'b0;
    n8013[78] = 1'b0;
    n8013[77] = 1'b0;
    n8013[76] = 1'b0;
    n8013[75] = 1'b0;
    n8013[74] = 1'b0;
    n8013[73] = 1'b0;
    n8013[72] = 1'b0;
    n8013[71] = 1'b0;
    n8013[70] = 1'b0;
    n8013[69] = 1'b0;
    n8013[68] = 1'b0;
    n8013[67] = 1'b0;
    n8013[66] = 1'b0;
    n8013[65] = 1'b0;
    n8013[64] = 1'b0;
    n8013[63] = 1'b0;
    n8013[62] = 1'b0;
    n8013[61] = 1'b0;
    n8013[60] = 1'b0;
    n8013[59] = 1'b0;
    n8013[58] = 1'b0;
    n8013[57] = 1'b0;
    n8013[56] = 1'b0;
    n8013[55] = 1'b0;
    n8013[54] = 1'b0;
    n8013[53] = 1'b0;
    n8013[52] = 1'b0;
    n8013[51] = 1'b0;
    n8013[50] = 1'b0;
    n8013[49] = 1'b0;
    n8013[48] = 1'b0;
    n8013[47] = 1'b0;
    n8013[46] = 1'b0;
    n8013[45] = 1'b0;
    n8013[44] = 1'b0;
    n8013[43] = 1'b0;
    n8013[42] = 1'b0;
    n8013[41] = 1'b0;
    n8013[40] = 1'b0;
    n8013[39] = 1'b0;
    n8013[38] = 1'b0;
    n8013[37] = 1'b0;
    n8013[36] = 1'b0;
    n8013[35] = 1'b0;
    n8013[34] = 1'b0;
    n8013[33] = 1'b0;
    n8013[32] = 1'b0;
    n8013[31] = 1'b0;
    n8013[30] = 1'b0;
    n8013[29] = 1'b0;
    n8013[28] = 1'b0;
    n8013[27] = 1'b0;
    n8013[26] = 1'b0;
    n8013[25] = 1'b0;
    n8013[24] = 1'b0;
    n8013[23] = 1'b0;
    n8013[22] = 1'b0;
    n8013[21] = 1'b0;
    n8013[20] = 1'b0;
    n8013[19] = 1'b0;
    n8013[18] = 1'b0;
    n8013[17] = 1'b0;
    n8013[16] = 1'b0;
    n8013[15] = 1'b0;
    n8013[14] = 1'b0;
    n8013[13] = 1'b0;
    n8013[12] = 1'b0;
    n8013[11] = 1'b0;
    n8013[10] = 1'b0;
    n8013[9] = 1'b0;
    n8013[8] = 1'b0;
    n8013[7] = 1'b0;
    n8013[6] = 1'b0;
    n8013[5] = 1'b0;
    n8013[4] = 1'b0;
    n8013[3] = 1'b0;
    n8013[2] = 1'b0;
    n8013[1] = 1'b0;
    n8013[0] = 1'b0;
    end
  assign n8014_data = n8013[n7727_o];
  /* decode1.vhdl:648:51  */
  /* decode1.vhdl:648:50  */
  reg [43:0] n8015[7:0] ; // memory
  initial begin
    n8015[7] = 44'b00000000000000000000110000000000000001110001;
    n8015[6] = 44'b00000000000000000000000010001000100000010001;
    n8015[5] = 44'b00000000000000000000000000000000000000000000;
    n8015[4] = 44'b00000000000000000000000000000000000000000000;
    n8015[3] = 44'b00010000000000000000010110001110011000111001;
    n8015[2] = 44'b00000000000000000000000000001110011101111001;
    n8015[1] = 44'b00000000000000000000000000000000000000000000;
    n8015[0] = 44'b00100000000000000000000000000000000011110001;
    end
  assign n8016_data = n8015[n7739_o];
  /* decode1.vhdl:650:44  */
  /* decode1.vhdl:650:43  */
  reg [43:0] n8017[15:0] ; // memory
  initial begin
    n8017[15] = 44'b00001000000000000000000100011100000110001001;
    n8017[14] = 44'b00001000000000000000000100011100000110001001;
    n8017[13] = 44'b00001000000000000000000100011100000110010001;
    n8017[12] = 44'b00001000000000000000000100011100000110010001;
    n8017[11] = 44'b00001000000000000000000100011100000110000001;
    n8017[10] = 44'b00001000000000000000000100011100000110000001;
    n8017[9] = 44'b00001000000000000000000100011100001110000001;
    n8017[8] = 44'b00001000000000000000000100011100001110000001;
    n8017[7] = 44'b00001000000000000000000100010001000110001001;
    n8017[6] = 44'b00001000000000000000000100010001000110010001;
    n8017[5] = 44'b00000000000000000000000000000000000000000000;
    n8017[4] = 44'b00000000000000000000000000000000000000000000;
    n8017[3] = 44'b00000000000000000000000000000000000000000000;
    n8017[2] = 44'b00000000000000000000000000000000000000000000;
    n8017[1] = 44'b00000000000000000000000000000000000000000000;
    n8017[0] = 44'b00000000000000000000000000000000000000000000;
    end
  assign n8018_data = n8017[n7804_o];
  /* decode1.vhdl:687:44  */
  /* decode1.vhdl:687:43  */
  reg [43:0] n8019[3:0] ; // memory
  initial begin
    n8019[3] = 44'b00000000000010000000000010001001010011111010;
    n8019[2] = 44'b11000000010010000000000010001001010011111010;
    n8019[1] = 44'b00000000001001100000000010001001010011111010;
    n8019[0] = 44'b00000000000000000000000000000000000000000000;
    end
  assign n8020_data = n8019[n7821_o];
  /* decode1.vhdl:696:44  */
  /* decode1.vhdl:696:43  */
  reg [43:0] n8021[31:0] ; // memory
  initial begin
    n8021[31] = 44'b00000000000000000000000000000000000000000000;
    n8021[30] = 44'b00000000000000000000000000000000000000000000;
    n8021[29] = 44'b00000000000000000000000000000000000000000000;
    n8021[28] = 44'b00000000000000000000000000000000000000000000;
    n8021[27] = 44'b00000000000000000000000000000000000000000000;
    n8021[26] = 44'b00000000000000000000000000000000000000000000;
    n8021[25] = 44'b00000000000000000000000000000000000000000000;
    n8021[24] = 44'b00000000000000000000000000000000000000000000;
    n8021[23] = 44'b00000000000000000000000000000000000000000000;
    n8021[22] = 44'b00000000000000000000000000000000000000000000;
    n8021[21] = 44'b00000000000000000000000000000000000000000000;
    n8021[20] = 44'b00000000000000000000000000000000000000000000;
    n8021[19] = 44'b00000000000000000000000000000000000000000000;
    n8021[18] = 44'b00000000000000000000000000000000000000000000;
    n8021[17] = 44'b00001001000000000000001000001111000011010111;
    n8021[16] = 44'b00000000000000000000000000000000000000000000;
    n8021[15] = 44'b00000000000000000000000000000000000000000000;
    n8021[14] = 44'b00000000000000000000000000000000000000000000;
    n8021[13] = 44'b00001001000000000000001000001111101011001111;
    n8021[12] = 44'b00000000000000000000000000000000000000000000;
    n8021[11] = 44'b00001001000000000000001000001111101011001111;
    n8021[10] = 44'b00001001000000000000001000001111101011001111;
    n8021[9] = 44'b00001001000000000000001000001111000011001111;
    n8021[8] = 44'b00000000000000000000000000000000000000000000;
    n8021[7] = 44'b00001001000000000000001000001111000011001111;
    n8021[6] = 44'b00001001000000000000001000110000101011001111;
    n8021[5] = 44'b00001001000000000000001000001111000011001111;
    n8021[4] = 44'b00000000000000000000000000000000000000000000;
    n8021[3] = 44'b00001001000000000000001000111111101011001111;
    n8021[2] = 44'b00001001000000000000001000111111101011001111;
    n8021[1] = 44'b00001001000000000000001000111111101011001111;
    n8021[0] = 44'b00001001000000000000001000111111101011001111;
    end
  assign n8022_data = n8021[n7830_o];
  /* decode1.vhdl:701:48  */
  /* decode1.vhdl:701:47  */
  reg [43:0] n8023[3:0] ; // memory
  initial begin
    n8023[3] = 44'b00000000000010000000000000011001010100000010;
    n8023[2] = 44'b00000000010010000000000100011001010100000010;
    n8023[1] = 44'b01000000000010000000000000011001010100000010;
    n8023[0] = 44'b00000000000000000000000000000000000000000000;
    end
  assign n8024_data = n8023[n7851_o];
  /* decode1.vhdl:708:44  */
  /* decode1.vhdl:708:43  */
  reg [43:0] n8025[511:0] ; // memory
  initial begin
    n8025[511] = 44'b00000000000000000000100000001111101011001111;
    n8025[510] = 44'b00000000000000000000100000001111101011001111;
    n8025[509] = 44'b00000000000000000000100000000000000011001111;
    n8025[508] = 44'b00000000000000000000000000000000000000000000;
    n8025[507] = 44'b00000000000000000000100000001111101011001111;
    n8025[506] = 44'b00000000000000000000100000001111000011001111;
    n8025[505] = 44'b00000000000000000000000000000000000000000000;
    n8025[504] = 44'b00000000000000000000000000000000000000000000;
    n8025[503] = 44'b00000000000000000000000000000000000000000000;
    n8025[502] = 44'b00000000000000000000000000000000000000000000;
    n8025[501] = 44'b00000000000000000000000000000000000000000000;
    n8025[500] = 44'b00000000000000000000000000000000000000000000;
    n8025[499] = 44'b00000000000000000000000000000000000000000000;
    n8025[498] = 44'b00000000000000000000000000000000000000000000;
    n8025[497] = 44'b00000000000000000000000000000000000000000000;
    n8025[496] = 44'b00000000000000000000000000000000000000000000;
    n8025[495] = 44'b00000000000000000000000000000000000000000000;
    n8025[494] = 44'b00000000000000000000000000000000000000000000;
    n8025[493] = 44'b00000000000000000000000000000000000000000000;
    n8025[492] = 44'b00000000000000000000000000000000000000000000;
    n8025[491] = 44'b00000000000000000000000000000000000000000000;
    n8025[490] = 44'b00000000000000000000000000000000000000000000;
    n8025[489] = 44'b00000000000000000000000000000000000000000000;
    n8025[488] = 44'b00000000000000000000000000000000000000000000;
    n8025[487] = 44'b00000000000000000000000000000000000000000000;
    n8025[486] = 44'b00000000000000000000000000000000000000000000;
    n8025[485] = 44'b00000000000000000000000000000000000000000000;
    n8025[484] = 44'b00000000000000000000000000000000000000000000;
    n8025[483] = 44'b00000000000000000000000000000000000000000000;
    n8025[482] = 44'b00000000000000000000000000000000000000000000;
    n8025[481] = 44'b00000000000000000000000000000000000000000000;
    n8025[480] = 44'b00000000000000000000000000000000000000000000;
    n8025[479] = 44'b00000000000000000000000000000000000000000000;
    n8025[478] = 44'b00000000000000000000000000000000000000000000;
    n8025[477] = 44'b00000000000000000000000000000000000000000000;
    n8025[476] = 44'b00000000000000000000000000000000000000000000;
    n8025[475] = 44'b00000000000000000000000000000000000000000000;
    n8025[474] = 44'b00000000000000000000000000000000000000000000;
    n8025[473] = 44'b00000000000000000000000000000000000000000000;
    n8025[472] = 44'b00000000000000000000000000000000000000000000;
    n8025[471] = 44'b00000000000000000000000000000000000000000000;
    n8025[470] = 44'b00000000000000000000000000000000000000000000;
    n8025[469] = 44'b00000000000000000000000000000000000000000000;
    n8025[468] = 44'b00000000000000000000000000000000000000000000;
    n8025[467] = 44'b00000000000000000000000000000000000000000000;
    n8025[466] = 44'b00000000000000000000000000000000000000000000;
    n8025[465] = 44'b00000000000000000000000000000000000000000000;
    n8025[464] = 44'b00000000000000000000000000000000000000000000;
    n8025[463] = 44'b00000000000000000000000000000000000000000000;
    n8025[462] = 44'b00000000000000000000000000000000000000000000;
    n8025[461] = 44'b00000000000000000000000000000000000000000000;
    n8025[460] = 44'b00000000000000000000000000000000000000000000;
    n8025[459] = 44'b00000000000000000000000000000000000000000000;
    n8025[458] = 44'b00000000000000000000000000000000000000000000;
    n8025[457] = 44'b00000000000000000000000000000000000000000000;
    n8025[456] = 44'b00000000000000000000000000000000000000000000;
    n8025[455] = 44'b00000000000000000000000000000000000000000000;
    n8025[454] = 44'b00000000000000000000000000000000000000000000;
    n8025[453] = 44'b00000000000000000000000000000000000000000000;
    n8025[452] = 44'b00000000000000000000000000000000000000000000;
    n8025[451] = 44'b00000000000000000000000000000000000000000000;
    n8025[450] = 44'b00000000000000000000000000000000000000000000;
    n8025[449] = 44'b00000000000000000000000000000000000000000000;
    n8025[448] = 44'b00000000000000000000000000000000000000000000;
    n8025[447] = 44'b00000000000000000000000000000000000000000000;
    n8025[446] = 44'b00000000000000000000000000000000000000000000;
    n8025[445] = 44'b00000000000000000000000000000000000000000000;
    n8025[444] = 44'b00000000000000000000000000000000000000000000;
    n8025[443] = 44'b00000000000000000000000000000000000000000000;
    n8025[442] = 44'b00000000000000000000000000000000000000000000;
    n8025[441] = 44'b00000000000000000000000000000000000000000000;
    n8025[440] = 44'b00000000000000000000000000000000000000000000;
    n8025[439] = 44'b00000000000000000000000000000000000000000000;
    n8025[438] = 44'b00000000000000000000000000000000000000000000;
    n8025[437] = 44'b00000000000000000000000000000000000000000000;
    n8025[436] = 44'b00000000000000000000000000000000000000000000;
    n8025[435] = 44'b00000000000000000000000000000000000000000000;
    n8025[434] = 44'b00000000000000000000000000000000000000000000;
    n8025[433] = 44'b00000000000000000000000000000000000000000000;
    n8025[432] = 44'b00000000000000000000000000000000000000000000;
    n8025[431] = 44'b00000000000000000000000000000000000000000000;
    n8025[430] = 44'b00000000000000000000000000000000000000000000;
    n8025[429] = 44'b00000000000000000000000000000000000000000000;
    n8025[428] = 44'b00000000000000000000000000000000000000000000;
    n8025[427] = 44'b00000000000000000000000000000000000000000000;
    n8025[426] = 44'b00000000000000000000000000000000000000000000;
    n8025[425] = 44'b00000000000000000000000000000000000000000000;
    n8025[424] = 44'b00000000000000000000000000000000000000000000;
    n8025[423] = 44'b00000000000000000000000000000000000000000000;
    n8025[422] = 44'b00000000000000000000000000000000000000000000;
    n8025[421] = 44'b00000000000000000000000000000000000000000000;
    n8025[420] = 44'b00000000000000000000000000000000000000000000;
    n8025[419] = 44'b00000000000000000000000000000000000000000000;
    n8025[418] = 44'b00000000000000000000000000000000000000000000;
    n8025[417] = 44'b00000000000000000000000000000000000000000000;
    n8025[416] = 44'b00000000000000000000000000000000000000000000;
    n8025[415] = 44'b00000000000000000000000000000000000000000000;
    n8025[414] = 44'b00000000000000000000000000000000000000000000;
    n8025[413] = 44'b00000000000000000000000000000000000000000000;
    n8025[412] = 44'b00000000000000000000000000000000000000000000;
    n8025[411] = 44'b00000000000000000000000000000000000000000000;
    n8025[410] = 44'b00000000000000000000000000000000000000000000;
    n8025[409] = 44'b00000000000000000000000000000000000000000000;
    n8025[408] = 44'b00000000000000000000000000000000000000000000;
    n8025[407] = 44'b00000000000000000000000000000000000000000000;
    n8025[406] = 44'b00000000000000000000000000000000000000000000;
    n8025[405] = 44'b00000000000000000000000000000000000000000000;
    n8025[404] = 44'b00000000000000000000000000000000000000000000;
    n8025[403] = 44'b00000000000000000000000000000000000000000000;
    n8025[402] = 44'b00000000000000000000000000000000000000000000;
    n8025[401] = 44'b00000000000000000000000000000000000000000000;
    n8025[400] = 44'b00000000000000000000000000000000000000000000;
    n8025[399] = 44'b00000000000000000000000000000000000000000000;
    n8025[398] = 44'b00000000000000000000000000000000000000000000;
    n8025[397] = 44'b00000000000000000000000000000000000000000000;
    n8025[396] = 44'b00000000000000000000000000000000000000000000;
    n8025[395] = 44'b00000000000000000000000000000000000000000000;
    n8025[394] = 44'b00000000000000000000000000000000000000000000;
    n8025[393] = 44'b00000000000000000000000000000000000000000000;
    n8025[392] = 44'b00000000000000000000000000000000000000000000;
    n8025[391] = 44'b00000000000000000000000000000000000000000000;
    n8025[390] = 44'b00000000000000000000000000000000000000000000;
    n8025[389] = 44'b00000000000000000000000000000000000000000000;
    n8025[388] = 44'b00000000000000000000000000000000000000000000;
    n8025[387] = 44'b00000000000000000000000000000000000000000000;
    n8025[386] = 44'b00000000000000000000000000000000000000000000;
    n8025[385] = 44'b00000000000000000000000000000000000000000000;
    n8025[384] = 44'b00000000000000000000000000000000000000000000;
    n8025[383] = 44'b00000000000000000000000000000000000000000000;
    n8025[382] = 44'b00000000000000000000000000000000000000000000;
    n8025[381] = 44'b00000000000000000000000000000000000000000000;
    n8025[380] = 44'b00000000000000000000000000000000000000000000;
    n8025[379] = 44'b00000000000000000000000000000000000000000000;
    n8025[378] = 44'b00000000000000000000000000000000000000000000;
    n8025[377] = 44'b00000000000000000000000000000000000000000000;
    n8025[376] = 44'b00000000000000000000000000000000000000000000;
    n8025[375] = 44'b00000000000000000000000000000000000000000000;
    n8025[374] = 44'b00000000000000000000000000000000000000000000;
    n8025[373] = 44'b00000000000000000000000000000000000000000000;
    n8025[372] = 44'b00000000000000000000000000000000000000000000;
    n8025[371] = 44'b00000000000000000000000000000000000000000000;
    n8025[370] = 44'b00000000000000000000000000000000000000000000;
    n8025[369] = 44'b00000000000000000000000000000000000000000000;
    n8025[368] = 44'b00000000000000000000000000000000000000000000;
    n8025[367] = 44'b00000000000000000000000000000000000000000000;
    n8025[366] = 44'b00000000000000000000000000000000000000000000;
    n8025[365] = 44'b00000000000000000000000000000000000000000000;
    n8025[364] = 44'b00000000000000000000000000000000000000000000;
    n8025[363] = 44'b00000000000000000000000000000000000000000000;
    n8025[362] = 44'b00000000000000000000000000000000000000000000;
    n8025[361] = 44'b00000000000000000000000000000000000000000000;
    n8025[360] = 44'b00000000000000000000000000000000000000000000;
    n8025[359] = 44'b00000000000000000000000000000000000000000000;
    n8025[358] = 44'b00000000000000000000000000000000000000000000;
    n8025[357] = 44'b00000000000000000000000000000000000000000000;
    n8025[356] = 44'b00000000000000000000000000000000000000000000;
    n8025[355] = 44'b00000000000000000000000000000000000000000000;
    n8025[354] = 44'b00000000000000000000000000000000000000000000;
    n8025[353] = 44'b00000000000000000000000000000000000000000000;
    n8025[352] = 44'b00000000000000000000000000000000000000000000;
    n8025[351] = 44'b00000000000000000000000000000000000000000000;
    n8025[350] = 44'b00000000000000000000000000000000000000000000;
    n8025[349] = 44'b00000000000000000000000000000000000000000000;
    n8025[348] = 44'b00000000000000000000000000000000000000000000;
    n8025[347] = 44'b00000000000000000000000000000000000000000000;
    n8025[346] = 44'b00000000000000000000000000000000000000000000;
    n8025[345] = 44'b00000000000000000000000000000000000000000000;
    n8025[344] = 44'b00000000000000000000000000000000000000000000;
    n8025[343] = 44'b00000000000000000000000000000000000000000000;
    n8025[342] = 44'b00000000000000000000000000000000000000000000;
    n8025[341] = 44'b00000000000000000000000000000000000000000000;
    n8025[340] = 44'b00000000000000000000000000000000000000000000;
    n8025[339] = 44'b00000000000000000000000000000000000000000000;
    n8025[338] = 44'b00000000000000000000000000000000000000000000;
    n8025[337] = 44'b00000000000000000000000000000000000000000000;
    n8025[336] = 44'b00000000000000000000000000000000000000000000;
    n8025[335] = 44'b00000000000000000000000000000000000000000000;
    n8025[334] = 44'b00000000000000000000000000000000000000000000;
    n8025[333] = 44'b00000000000000000000000000000000000000000000;
    n8025[332] = 44'b00000000000000000000000000000000000000000000;
    n8025[331] = 44'b00000000000000000000000000000000000000000000;
    n8025[330] = 44'b00000000000000000000000000000000000000000000;
    n8025[329] = 44'b00000000000000000000000000000000000000000000;
    n8025[328] = 44'b00000000000000000000000000000000000000000000;
    n8025[327] = 44'b00000000000000000000000000000000000000000000;
    n8025[326] = 44'b00000000000000000000000000000000000000000000;
    n8025[325] = 44'b00000000000000000000000000000000000000000000;
    n8025[324] = 44'b00000000000000000000000000000000000000000000;
    n8025[323] = 44'b00000000000000000000000000000000000000000000;
    n8025[322] = 44'b00000000000000000000000000000000000000000000;
    n8025[321] = 44'b00000000000000000000000000000000000000000000;
    n8025[320] = 44'b00000000000000000000000000000000000000000000;
    n8025[319] = 44'b00000000000000000000000000000000000000000000;
    n8025[318] = 44'b00001000000000000000000000000000000011001111;
    n8025[317] = 44'b00001000000000000000000000000000000011001111;
    n8025[316] = 44'b00000000000000000000000000000000000000000000;
    n8025[315] = 44'b00001000000000000000000000000000000011001111;
    n8025[314] = 44'b00000000000000000000000000000000000000000000;
    n8025[313] = 44'b00000000000000000000000000000000000000000000;
    n8025[312] = 44'b00000000000000000000000000000000000000000000;
    n8025[311] = 44'b00000000000000000000000000000000000000000000;
    n8025[310] = 44'b00000000000000000000000000000000000000000000;
    n8025[309] = 44'b00000000000000000000000000000000000000000000;
    n8025[308] = 44'b00000000000000000000000000000000000000000000;
    n8025[307] = 44'b00000000000000000000000000000000000000000000;
    n8025[306] = 44'b00000000000000000000000000000000000000000000;
    n8025[305] = 44'b00000000000000000000000000000000000000000000;
    n8025[304] = 44'b00000000000000000000000000000000000000000000;
    n8025[303] = 44'b00000000000000000000000000000000000000000000;
    n8025[302] = 44'b00000000000000000000000000000000000000000000;
    n8025[301] = 44'b00000000000000000000000000000000000000000000;
    n8025[300] = 44'b00000000000000000000000000000000000000000000;
    n8025[299] = 44'b00000000000000000000000000000000000000000000;
    n8025[298] = 44'b00000000000000000000000000000000000000000000;
    n8025[297] = 44'b00000000000000000000000000000000000000000000;
    n8025[296] = 44'b00000000000000000000000000000000000000000000;
    n8025[295] = 44'b00000000000000000000000000000000000000000000;
    n8025[294] = 44'b00000000000000000000000000000000000000000000;
    n8025[293] = 44'b00000000000000000000001000001111101011010111;
    n8025[292] = 44'b00000000000000000000000000000000000000000000;
    n8025[291] = 44'b00000000000000000000000000000000000000000000;
    n8025[290] = 44'b00000000000000000000000000000000000000000000;
    n8025[289] = 44'b00000000000000000000001000001111101011010111;
    n8025[288] = 44'b00000000000000000000000000000000000000000000;
    n8025[287] = 44'b00000000000000000000000000000000000000000000;
    n8025[286] = 44'b00000000000000000000000000000000000000000000;
    n8025[285] = 44'b00000000000000000000000000000000000000000000;
    n8025[284] = 44'b00000000000000000000000000000000000000000000;
    n8025[283] = 44'b00000000000000000000000000000000000000000000;
    n8025[282] = 44'b00000000000000000000000000000000000000000000;
    n8025[281] = 44'b00000000000000000000000000000000000000000000;
    n8025[280] = 44'b00000000000000000000000000000000000000000000;
    n8025[279] = 44'b00000000000000000000000000000000000000000000;
    n8025[278] = 44'b00000000000000000000000000000000000000000000;
    n8025[277] = 44'b00000000000000000000000000000000000000000000;
    n8025[276] = 44'b00000000000000000000000000000000000000000000;
    n8025[275] = 44'b00000000000000000000000000000000000000000000;
    n8025[274] = 44'b00000000000000000000000000000000000000000000;
    n8025[273] = 44'b00000000000000000000000000000000000000000000;
    n8025[272] = 44'b00000000000000000000000000000000000000000000;
    n8025[271] = 44'b00000000000000000000000000000000000000000000;
    n8025[270] = 44'b00000000000000000000000000000000000000000000;
    n8025[269] = 44'b00001000000000000000001000001111000011010111;
    n8025[268] = 44'b00000000000000000000000000000000000000000000;
    n8025[267] = 44'b00000000000000000000000000000000000000000000;
    n8025[266] = 44'b00000000000000000000000000000000000000000000;
    n8025[265] = 44'b00001000000000000000000000001111000011010111;
    n8025[264] = 44'b00000000000000000000000000000000000000000000;
    n8025[263] = 44'b00000000000000000000000000000000000000000000;
    n8025[262] = 44'b00000000000000000000000000000000000000000000;
    n8025[261] = 44'b00000000000000000000000000000000000000000000;
    n8025[260] = 44'b00000000000000000000000000000000000000000000;
    n8025[259] = 44'b00000000000000000000000000000000000000000000;
    n8025[258] = 44'b00000000000000000000000000000000000000000000;
    n8025[257] = 44'b00000000000000000000000000000000000000000000;
    n8025[256] = 44'b00000000000000000000000000000000000000000000;
    n8025[255] = 44'b00001000000000000000001000001111101011001111;
    n8025[254] = 44'b00001000000000000000001000001111000011001111;
    n8025[253] = 44'b00001000000000000000001000001111000011001111;
    n8025[252] = 44'b00000000000000000000000000000000000000000000;
    n8025[251] = 44'b00001000000000000000001000001111000011001111;
    n8025[250] = 44'b00000000000000000000000000000000000000000000;
    n8025[249] = 44'b00000000000000000000000000000000000000000000;
    n8025[248] = 44'b00000000000000000000000000000000000000000000;
    n8025[247] = 44'b00001000000000000000001000001111000011001111;
    n8025[246] = 44'b00000000000000000000000000000000000000000000;
    n8025[245] = 44'b00000000000000000000000000000000000000000000;
    n8025[244] = 44'b00000000000000000000000000000000000000000000;
    n8025[243] = 44'b00001000000000000000001000001111000011001111;
    n8025[242] = 44'b00001000000000000000001000001111000011001111;
    n8025[241] = 44'b00001000000000000000001000001111000011001111;
    n8025[240] = 44'b00001000000000000000001000001111000011001111;
    n8025[239] = 44'b00000000000000000000000000000000000000000000;
    n8025[238] = 44'b00000000000000000000000000000000000000000000;
    n8025[237] = 44'b00000000000000000000000000000000000000000000;
    n8025[236] = 44'b00000000000000000000000000000000000000000000;
    n8025[235] = 44'b00000000000000000000000000000000000000000000;
    n8025[234] = 44'b00000000000000000000000000000000000000000000;
    n8025[233] = 44'b00000000000000000000000000000000000000000000;
    n8025[232] = 44'b00000000000000000000000000000000000000000000;
    n8025[231] = 44'b00000000000000000000000000000000000000000000;
    n8025[230] = 44'b00000000000000000000000000000000000000000000;
    n8025[229] = 44'b00000000000000000000000000000000000000000000;
    n8025[228] = 44'b00000000000000000000000000000000000000000000;
    n8025[227] = 44'b00000000000000000000000000000000000000000000;
    n8025[226] = 44'b00000000000000000000000000000000000000000000;
    n8025[225] = 44'b00000000000000000000000000000000000000000000;
    n8025[224] = 44'b00000000000000000000000000000000000000000000;
    n8025[223] = 44'b00000000000000000000000000000000000000000000;
    n8025[222] = 44'b00000000000000000000000000000000000000000000;
    n8025[221] = 44'b00000000000000000000000000000000000000000000;
    n8025[220] = 44'b00000000000000000000000000000000000000000000;
    n8025[219] = 44'b00000000000000000000000000000000000000000000;
    n8025[218] = 44'b00000000000000000000000000000000000000000000;
    n8025[217] = 44'b00000000000000000000000000000000000000000000;
    n8025[216] = 44'b00000000000000000000000000000000000000000000;
    n8025[215] = 44'b00000000000000000000000000000000000000000000;
    n8025[214] = 44'b00000000000000000000000000000000000000000000;
    n8025[213] = 44'b00000000000000000000000000000000000000000000;
    n8025[212] = 44'b00000000000000000000000000000000000000000000;
    n8025[211] = 44'b00000000000000000000000000000000000000000000;
    n8025[210] = 44'b00000000000000000000000000000000000000000000;
    n8025[209] = 44'b00000000000000000000000000000000000000000000;
    n8025[208] = 44'b00000000000000000000000000000000000000000000;
    n8025[207] = 44'b00000000000000000000000000000000000000000000;
    n8025[206] = 44'b00000000000000000000000000000000000000000000;
    n8025[205] = 44'b00000000000000000000000000000000000000000000;
    n8025[204] = 44'b00000000000000000000000000000000000000000000;
    n8025[203] = 44'b00000000000000000000000000000000000000000000;
    n8025[202] = 44'b00000000000000000000000000000000000000000000;
    n8025[201] = 44'b00000000000000000000000000000000000000000000;
    n8025[200] = 44'b00000000000000000000000000000000000000000000;
    n8025[199] = 44'b00000000000000000000000000000000000000000000;
    n8025[198] = 44'b00000000000000000000000000000000000000000000;
    n8025[197] = 44'b00000000000000000000000000000000000000000000;
    n8025[196] = 44'b00000000000000000000000000000000000000000000;
    n8025[195] = 44'b00000000000000000000000000000000000000000000;
    n8025[194] = 44'b00000000000000000000000000000000000000000000;
    n8025[193] = 44'b00000000000000000000000000000000000000000000;
    n8025[192] = 44'b00000000000000000000000000000000000000000000;
    n8025[191] = 44'b00000000000000000000000000000000000000000000;
    n8025[190] = 44'b00000000000000000000000000000000000000000000;
    n8025[189] = 44'b00000000000000000000000000000000000000000000;
    n8025[188] = 44'b00000000000000000000000000000000000000000000;
    n8025[187] = 44'b00000000000000000000000000000000000000000000;
    n8025[186] = 44'b00000000000000000000000000000000000000000000;
    n8025[185] = 44'b00000000000000000000000000000000000000000000;
    n8025[184] = 44'b00000000000000000000000000000000000000000000;
    n8025[183] = 44'b00000000000000000000000000000000000000000000;
    n8025[182] = 44'b00000000000000000000000000000000000000000000;
    n8025[181] = 44'b00000000000000000000000000000000000000000000;
    n8025[180] = 44'b00000000000000000000000000000000000000000000;
    n8025[179] = 44'b00000000000000000000000000000000000000000000;
    n8025[178] = 44'b00000000000000000000000000000000000000000000;
    n8025[177] = 44'b00000000000000000000000000000000000000000000;
    n8025[176] = 44'b00000000000000000000000000000000000000000000;
    n8025[175] = 44'b00000000000000000000000000000000000000000000;
    n8025[174] = 44'b00000000000000000000000000000000000000000000;
    n8025[173] = 44'b00000000000000000000000000000000000000000000;
    n8025[172] = 44'b00000000000000000000000000000000000000000000;
    n8025[171] = 44'b00000000000000000000000000000000000000000000;
    n8025[170] = 44'b00000000000000000000000000000000000000000000;
    n8025[169] = 44'b00000000000000000000000000000000000000000000;
    n8025[168] = 44'b00000000000000000000000000000000000000000000;
    n8025[167] = 44'b00000000000000000000000000000000000000000000;
    n8025[166] = 44'b00000000000000000000000000000000000000000000;
    n8025[165] = 44'b00000000000000000000000000000000000000000000;
    n8025[164] = 44'b00000000000000000000000000000000000000000000;
    n8025[163] = 44'b00000000000000000000000000000000000000000000;
    n8025[162] = 44'b00000000000000000000000000000000000000000000;
    n8025[161] = 44'b00000000000000000000000000000000000000000000;
    n8025[160] = 44'b00000000000000000000000000000000000000000000;
    n8025[159] = 44'b00000000000000000000000000000000000000000000;
    n8025[158] = 44'b00000000000000000000000000000000000000000000;
    n8025[157] = 44'b00000000000000000000000000000000000000000000;
    n8025[156] = 44'b00000000000000000000000000000000000000000000;
    n8025[155] = 44'b00000000000000000000000000000000000000000000;
    n8025[154] = 44'b00000000000000000000000000000000000000000000;
    n8025[153] = 44'b00000000000000000000000000000000000000000000;
    n8025[152] = 44'b00000000000000000000000000000000000000000000;
    n8025[151] = 44'b00000000000000000000000000000000000000000000;
    n8025[150] = 44'b00000000000000000000000000000000000000000000;
    n8025[149] = 44'b00000000000000000000000000000000000000000000;
    n8025[148] = 44'b00000000000000000000000000000000000000000000;
    n8025[147] = 44'b00000000000000000000000000000000000000000000;
    n8025[146] = 44'b00000000000000000000000000000000000000000000;
    n8025[145] = 44'b00000000000000000000000000000000000000000000;
    n8025[144] = 44'b00000000000000000000000000000000000000000000;
    n8025[143] = 44'b00000000000000000000000000000000000000000000;
    n8025[142] = 44'b00000000000000000000000000000000000000000000;
    n8025[141] = 44'b00000000000000000000000000000000000000000000;
    n8025[140] = 44'b00000000000000000000000000000000000000000000;
    n8025[139] = 44'b00000000000000000000000000000000000000000000;
    n8025[138] = 44'b00000000000000000000000000000000000000000000;
    n8025[137] = 44'b00000000000000000000000000000000000000000000;
    n8025[136] = 44'b00000000000000000000000000000000000000000000;
    n8025[135] = 44'b00000000000000000000000000000000000000000000;
    n8025[134] = 44'b00000000000000000000000000000000000000000000;
    n8025[133] = 44'b00000000000000000000000000000000000000000000;
    n8025[132] = 44'b00000000000000000000000000000000000000000000;
    n8025[131] = 44'b00000000000000000000000000000000000000000000;
    n8025[130] = 44'b00000000000000000000000000000000000000000000;
    n8025[129] = 44'b00000000000000000000000000000000000000000000;
    n8025[128] = 44'b00000000000000000000000000000000000000000000;
    n8025[127] = 44'b00001001000000000000001000001111000011001111;
    n8025[126] = 44'b00000000000000000000000000000000000000000000;
    n8025[125] = 44'b00000000000000000000000000000000000000000000;
    n8025[124] = 44'b00000000000000000000000000000000000000000000;
    n8025[123] = 44'b00000000000000000000000000000000000000000000;
    n8025[122] = 44'b00000000000000000000000000000000000000000000;
    n8025[121] = 44'b00000000000000000000000000000000000000000000;
    n8025[120] = 44'b00000000000000000000000000000000000000000000;
    n8025[119] = 44'b00000000000000000000000000000000000000000000;
    n8025[118] = 44'b00000000000000000000000000000000000000000000;
    n8025[117] = 44'b00000000000000000000000000000000000000000000;
    n8025[116] = 44'b00000000000000000000000000000000000000000000;
    n8025[115] = 44'b00000000000000000000000000000000000000000000;
    n8025[114] = 44'b00000000000000000000000000000000000000000000;
    n8025[113] = 44'b00000000000000000000000000000000000000000000;
    n8025[112] = 44'b00000000000000000000000000000000000000000000;
    n8025[111] = 44'b00000000000000000000000000000000000000000000;
    n8025[110] = 44'b00000000000000000000000000000000000000000000;
    n8025[109] = 44'b00000000000000000000000000000000000000000000;
    n8025[108] = 44'b00000000000000000000000000000000000000000000;
    n8025[107] = 44'b00000000000000000000000000000000000000000000;
    n8025[106] = 44'b00000000000000000000000000000000000000000000;
    n8025[105] = 44'b00000000000000000000000000000000000000000000;
    n8025[104] = 44'b00000000000000000000000000000000000000000000;
    n8025[103] = 44'b00000000000000000000000000000000000000000000;
    n8025[102] = 44'b00000000000000000000000000000000000000000000;
    n8025[101] = 44'b00000000000000000000000000000000000000000000;
    n8025[100] = 44'b00000000000000000000000000000000000000000000;
    n8025[99] = 44'b00000000000000000000000000000000000000000000;
    n8025[98] = 44'b00000000000000000000000000000000000000000000;
    n8025[97] = 44'b00000000000000000000000000000000000000000000;
    n8025[96] = 44'b00000000000000000000000000000000000000000000;
    n8025[95] = 44'b00000000000000000000000000000000000000000000;
    n8025[94] = 44'b00000000000000000000000000000000000000000000;
    n8025[93] = 44'b00000000000000000000000000000000000000000000;
    n8025[92] = 44'b00000000000000000000000000000000000000000000;
    n8025[91] = 44'b00000000000000000000000000000000000000000000;
    n8025[90] = 44'b00000000000000000000000000000000000000000000;
    n8025[89] = 44'b00000000000000000000000000000000000000000000;
    n8025[88] = 44'b00000000000000000000000000000000000000000000;
    n8025[87] = 44'b00000000000000000000000000000000000000000000;
    n8025[86] = 44'b00000000000000000000000000000000000000000000;
    n8025[85] = 44'b00000000000000000000000000000000000000000000;
    n8025[84] = 44'b00000000000000000000000000000000000000000000;
    n8025[83] = 44'b00000000000000000000000000000000000000000000;
    n8025[82] = 44'b00000000000000000000000000000000000000000000;
    n8025[81] = 44'b00000000000000000000000000000000000000000000;
    n8025[80] = 44'b00000000000000000000000000000000000000000000;
    n8025[79] = 44'b00000000000000000000000000000000000000000000;
    n8025[78] = 44'b00000000000000000000000000000000000000000000;
    n8025[77] = 44'b00000000000000000000000000000000000000000000;
    n8025[76] = 44'b00000000000000000000000000000000000000000000;
    n8025[75] = 44'b00000000000000000000000000000000000000000000;
    n8025[74] = 44'b00000000000000000000000000000000000000000000;
    n8025[73] = 44'b00000000000000000000000000000000000000000000;
    n8025[72] = 44'b00000000000000000000000000000000000000000000;
    n8025[71] = 44'b00000000000000000000000000000000000000000000;
    n8025[70] = 44'b00000000000000000000000000000000000000000000;
    n8025[69] = 44'b00000000000000000000000000000000000000000000;
    n8025[68] = 44'b00000000000000000000000000000000000000000000;
    n8025[67] = 44'b00000000000000000000000000000000000000000000;
    n8025[66] = 44'b00000000000000000000000000000000000000000000;
    n8025[65] = 44'b00000000000000000000000000000000000000000000;
    n8025[64] = 44'b00000000000000000000000000000000000000000000;
    n8025[63] = 44'b00001000000000000000001000001111000011001111;
    n8025[62] = 44'b00000000000000000000000000000000000000000000;
    n8025[61] = 44'b00000000000000000000000000000000000000000000;
    n8025[60] = 44'b00000000000000000000000000000000000000000000;
    n8025[59] = 44'b00001000000000000000001000001111000011001111;
    n8025[58] = 44'b00000000000000000000000000000000000000000000;
    n8025[57] = 44'b00000000000000000000000000000000000000000000;
    n8025[56] = 44'b00000000000000000000000000000000000000000000;
    n8025[55] = 44'b00000000000000000000000000000000000000000000;
    n8025[54] = 44'b00000000000000000000000000000000000000000000;
    n8025[53] = 44'b00000000000000000000000000000000000000000000;
    n8025[52] = 44'b00000000000000000000000000000000000000000000;
    n8025[51] = 44'b00000000000000000000000000000000000000000000;
    n8025[50] = 44'b00000000000000000000000000000000000000000000;
    n8025[49] = 44'b00000000000000000000000000000000000000000000;
    n8025[48] = 44'b00000000000000000000000000000000000000000000;
    n8025[47] = 44'b00000000000000000000000000000000000000000000;
    n8025[46] = 44'b00000000000000000000000000000000000000000000;
    n8025[45] = 44'b00000000000000000000000000000000000000000000;
    n8025[44] = 44'b00000000000000000000000000000000000000000000;
    n8025[43] = 44'b00000000000000000000000000000000000000000000;
    n8025[42] = 44'b00000000000000000000000000000000000000000000;
    n8025[41] = 44'b00000000000000000000000000000000000000000000;
    n8025[40] = 44'b00000000000000000000000000000000000000000000;
    n8025[39] = 44'b00000000000000000000000000000000000000000000;
    n8025[38] = 44'b00001000000000000000001000001111000011001111;
    n8025[37] = 44'b00001000000000000000001000001111000011010111;
    n8025[36] = 44'b00000000000000000000000000000000000000000000;
    n8025[35] = 44'b00000000000000000000000000000000000000000000;
    n8025[34] = 44'b00001000000000000000001000001111000011001111;
    n8025[33] = 44'b00001000000000000000001000001111000011010111;
    n8025[32] = 44'b00000000000000000000000000000000000000000000;
    n8025[31] = 44'b00001000000000000000001000001111000011001111;
    n8025[30] = 44'b00000000000000000000000000000000000000000000;
    n8025[29] = 44'b00000000000000000000000000000000000000000000;
    n8025[28] = 44'b00000000000000000000000000000000000000000000;
    n8025[27] = 44'b00001000000000000000001000001111000011001111;
    n8025[26] = 44'b00000000000000000000000000000000000000000000;
    n8025[25] = 44'b00000000000000000000000000000000000000000000;
    n8025[24] = 44'b00000000000000000000000000000000000000000000;
    n8025[23] = 44'b00000000000000000000000000000000000000000000;
    n8025[22] = 44'b00000000000000000000000000000000000000000000;
    n8025[21] = 44'b00000000000000000000000000000000000000000000;
    n8025[20] = 44'b00000000000000000000000000000000000000000000;
    n8025[19] = 44'b00000000000000000000000000000000000000000000;
    n8025[18] = 44'b00000000000000000000000000000000000000000000;
    n8025[17] = 44'b00000000000000000000000000000000000000000000;
    n8025[16] = 44'b00000000000000000000000000000000000000000000;
    n8025[15] = 44'b00000000000000000000000000000000000000000000;
    n8025[14] = 44'b00000000000000000000000000000000000000000000;
    n8025[13] = 44'b00000000000000000000000000000000000000000000;
    n8025[12] = 44'b00000000000000000000000000000000000000000000;
    n8025[11] = 44'b00000000000000000000000000000000000000000000;
    n8025[10] = 44'b00000000000000000000000000000000000000000000;
    n8025[9] = 44'b00000000000000000000000000000000000000000000;
    n8025[8] = 44'b00000000000000000000000000000000000000000000;
    n8025[7] = 44'b00000000000000000000000000000000000000000000;
    n8025[6] = 44'b00001000000000000000001000001111000011001111;
    n8025[5] = 44'b00000000000000000000000000000000000000000000;
    n8025[4] = 44'b00000000000000000000000000000000000000000000;
    n8025[3] = 44'b00000000000000000000000000000000000000000000;
    n8025[2] = 44'b00001000000000000000001000001111000011001111;
    n8025[1] = 44'b00000000000000000000000000000000000000000000;
    n8025[0] = 44'b00000000000000000000000000000000000000000000;
    end
  assign n8026_data = n8025[n7864_o];
  /* decode1.vhdl:714:53  */
  /* decode1.vhdl:714:52  */
  reg [43:0] n8027[16:0] ; // memory
  initial begin
    n8027[16] = 44'b00000000000000000000000000000000000000000000;
    n8027[15] = 44'b00000000000000000000000000000000000000000000;
    n8027[14] = 44'b00001000000000000000001000001111101011001111;
    n8027[13] = 44'b00000000000000000000000000000000000000000000;
    n8027[12] = 44'b00001000000000000000001000001111101011001111;
    n8027[11] = 44'b00001000000000000000001000001111101011001111;
    n8027[10] = 44'b00001000000000000000001000001111000011001111;
    n8027[9] = 44'b00001000000000000000001000111111101011001111;
    n8027[8] = 44'b00001000000000000000001000001111000011001111;
    n8027[7] = 44'b00001000000000000000001000110000101011001111;
    n8027[6] = 44'b00001000000000000000001000001111000011001111;
    n8027[5] = 44'b00000000000000000000000000000000000000000000;
    n8027[4] = 44'b00001000000000000000001000111111101011001111;
    n8027[3] = 44'b00001000000000000000001000111111101011001111;
    n8027[2] = 44'b00001000000000000000001000111111101011001111;
    n8027[1] = 44'b00001000000000000000001000111111101011001111;
    n8027[0] = 44'b00000000000000000000000000000000000000000000;
    end
  assign n8028_data = n8027[n7872_o];
  /* decode1.vhdl:716:53  */
endmodule

module icache_64_8_4_1_4_12_0_5ba93c9db0cff93f52b521d7420e43f6eda2784f
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  clk,
   input  rst,
   input  i_in_req,
   input  i_in_virt_mode,
   input  i_in_priv_mode,
   input  i_in_big_endian,
   input  i_in_stop_mark,
   input  i_in_predicted,
   input  i_in_pred_ntaken,
   input  [63:0] i_in_nia,
   input  m_in_tlbld,
   input  m_in_tlbie,
   input  m_in_doall,
   input  [63:0] m_in_addr,
   input  [63:0] m_in_pte,
   input  stall_in,
   input  flush_in,
   input  inval_in,
   input  [63:0] wishbone_in_dat,
   input  wishbone_in_ack,
   input  wishbone_in_stall,
   input  [28:0] wb_snoop_in_adr,
   input  [63:0] wb_snoop_in_dat,
   input  [7:0] wb_snoop_in_sel,
   input  wb_snoop_in_cyc,
   input  wb_snoop_in_stb,
   input  wb_snoop_in_we,
   output i_out_valid,
   output i_out_stop_mark,
   output i_out_fetch_failed,
   output [63:0] i_out_nia,
   output [31:0] i_out_insn,
   output i_out_big_endian,
   output i_out_next_predicted,
   output i_out_next_pred_ntaken,
   output stall_out,
   output [28:0] wishbone_out_adr,
   output [63:0] wishbone_out_dat,
   output [7:0] wishbone_out_sel,
   output wishbone_out_cyc,
   output wishbone_out_stb,
   output wishbone_out_we,
   output events_icache_miss,
   output events_itlb_miss_resolved,
   output [53:0] log_out);
  wire [70:0] n6287_o;
  wire n6289_o;
  wire n6290_o;
  wire n6291_o;
  wire [63:0] n6292_o;
  wire [31:0] n6293_o;
  wire n6294_o;
  wire n6295_o;
  wire n6296_o;
  wire [130:0] n6297_o;
  wire [28:0] n6300_o;
  wire [63:0] n6301_o;
  wire [7:0] n6302_o;
  wire n6303_o;
  wire n6304_o;
  wire n6305_o;
  wire [65:0] n6306_o;
  wire [103:0] n6307_o;
  wire n6309_o;
  wire n6310_o;
  wire [195:0] cache_tags;
  wire [3:0] cache_valids;
  wire [3:0] itlb_valids;
  wire eaa_priv;
  wire [241:0] r;
  wire [1:0] req_index;
  wire [4:0] req_row;
  wire [48:0] req_tag;
  wire req_is_hit;
  wire req_is_miss;
  wire [55:0] req_raddr;
  wire [1:0] tlb_req_index;
  wire [55:0] real_addr;
  wire ra_valid;
  wire priv_fault;
  wire access_ok;
  wire [63:0] cache_out;
  wire snoop_valid;
  wire [1:0] snoop_index;
  wire snoop_hits;
  wire rams_n1_do_read;
  wire rams_n1_do_write;
  wire [4:0] rams_n1_rd_addr;
  wire [4:0] rams_n1_wr_addr;
  wire [63:0] rams_n1_dout;
  wire [7:0] rams_n1_wr_sel;
  wire [63:0] rams_n1_wr_dat;
  wire [63:0] rams_n1_way_rd_data;
  wire n6320_o;
  wire n6321_o;
  wire [63:0] n6322_o;
  wire [7:0] n6323_o;
  wire [7:0] n6324_o;
  wire [7:0] n6325_o;
  wire [7:0] n6326_o;
  wire [7:0] n6327_o;
  wire [7:0] n6328_o;
  wire [7:0] n6329_o;
  wire [7:0] n6330_o;
  wire [63:0] n6331_o;
  wire [63:0] n6332_o;
  wire n6335_o;
  wire n6336_o;
  wire n6338_o;
  wire n6341_o;
  wire [4:0] n6344_o;
  wire [7:0] n6347_o;
  wire [63:0] n6352_o;
  wire [1:0] n6358_o;
  wire [1:0] n6359_o;
  wire [1:0] n6360_o;
  wire [1:0] n6361_o;
  wire [1:0] n6362_o;
  wire n6373_o;
  wire [43:0] n6374_o;
  wire [11:0] n6375_o;
  wire [55:0] n6376_o;
  wire [49:0] n6377_o;
  wire n6378_o;
  wire [1:0] n6380_o;
  wire n6384_o;
  wire n6385_o;
  wire [63:0] n6387_o;
  wire [55:0] n6392_o;
  wire n6394_o;
  wire [55:0] n6395_o;
  wire n6397_o;
  wire n6398_o;
  wire n6399_o;
  wire n6400_o;
  wire n6401_o;
  wire n6402_o;
  wire [63:0] n6408_o;
  wire [1:0] n6414_o;
  wire [1:0] n6415_o;
  wire [1:0] n6416_o;
  wire [1:0] n6417_o;
  wire [1:0] n6418_o;
  wire n6421_o;
  wire n6422_o;
  wire n6423_o;
  wire n6424_o;
  wire n6429_o;
  wire [1:0] n6431_o;
  wire n6435_o;
  wire [49:0] n6439_o;
  wire [63:0] n6444_o;
  wire [1:0] n6447_o;
  wire [3:0] n6451_o;
  wire [3:0] n6454_o;
  wire [3:0] n6457_o;
  wire [3:0] n6458_o;
  wire [63:0] n6475_o;
  wire [1:0] n6480_o;
  wire [63:0] n6483_o;
  wire [4:0] n6488_o;
  wire n6491_o;
  wire [47:0] n6496_o;
  wire [48:0] n6497_o;
  wire [52:0] n6498_o;
  wire [55:0] n6500_o;
  wire n6501_o;
  wire [1:0] n6503_o;
  wire [1:0] n6506_o;
  wire n6508_o;
  wire [31:0] n6509_o;
  wire [1:0] n6510_o;
  wire [31:0] n6511_o;
  wire n6512_o;
  wire n6513_o;
  wire n6515_o;
  wire [31:0] n6516_o;
  wire [2:0] n6517_o;
  wire [2:0] n6520_o;
  wire n6523_o;
  wire n6524_o;
  wire n6525_o;
  wire [1:0] n6528_o;
  wire n6535_o;
  wire n6538_o;
  wire n6540_o;
  wire n6542_o;
  wire n6543_o;
  wire n6544_o;
  wire n6545_o;
  wire n6546_o;
  wire n6547_o;
  wire n6548_o;
  wire n6550_o;
  wire n6552_o;
  wire [63:0] n6563_o;
  wire n6569_o;
  wire n6582_o;
  wire [63:0] n6583_o;
  wire n6584_o;
  wire n6585_o;
  wire n6586_o;
  wire n6587_o;
  wire n6588_o;
  wire n6589_o;
  wire n6590_o;
  wire [103:0] n6591_o;
  wire n6597_o;
  wire n6599_o;
  wire n6600_o;
  wire n6601_o;
  wire n6602_o;
  wire n6603_o;
  wire [63:0] n6604_o;
  wire n6605_o;
  wire [64:0] n6606_o;
  wire [64:0] n6607_o;
  wire [64:0] n6608_o;
  wire n6609_o;
  wire n6610_o;
  wire [66:0] n6611_o;
  wire n6634_o;
  wire n6635_o;
  wire n6636_o;
  wire n6637_o;
  wire n6638_o;
  wire [28:0] n6641_o;
  localparam [63:0] n6647_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] n6648_o;
  wire [2:0] n6649_o;
  wire [63:0] n6650_o;
  wire [55:0] n6655_o;
  wire [1:0] n6661_o;
  wire [1:0] n6668_o;
  wire [1:0] n6671_o;
  wire [47:0] n6679_o;
  wire [48:0] n6681_o;
  wire [47:0] n6688_o;
  wire [48:0] n6689_o;
  wire n6690_o;
  wire n6693_o;
  wire n6700_o;
  wire [1:0] n6702_o;
  wire [3:0] n6706_o;
  wire [3:0] n6707_o;
  wire [3:0] n6708_o;
  wire n6709_o;
  wire n6710_o;
  wire [1:0] n6711_o;
  wire [4:0] n6726_o;
  wire [4:0] n6735_o;
  wire [2:0] n6744_o;
  wire [2:0] n6746_o;
  wire [28:0] n6752_o;
  wire [30:0] n6756_o;
  wire [1:0] n6757_o;
  wire [59:0] n6758_o;
  wire [30:0] n6759_o;
  wire [30:0] n6760_o;
  wire [1:0] n6761_o;
  wire [1:0] n6762_o;
  wire [55:0] n6763_o;
  wire [2:0] n6764_o;
  wire [59:0] n6765_o;
  wire [59:0] n6766_o;
  wire n6769_o;
  wire [1:0] n6770_o;
  wire n6772_o;
  wire [1:0] n6774_o;
  wire [48:0] n6784_o;
  wire [1:0] n6787_o;
  wire [1:0] n6789_o;
  wire [195:0] n6793_o;
  wire [3:0] n6794_o;
  wire [1:0] n6795_o;
  wire [1:0] n6796_o;
  wire n6798_o;
  wire n6799_o;
  wire [103:0] n6800_o;
  wire n6801_o;
  wire n6802_o;
  wire [103:0] n6804_o;
  wire [28:0] n6805_o;
  wire [2:0] n6806_o;
  wire [2:0] n6811_o;
  wire n6812_o;
  wire n6814_o;
  wire n6815_o;
  wire [103:0] n6817_o;
  wire [28:0] n6818_o;
  wire [2:0] n6825_o;
  wire [2:0] n6828_o;
  wire [25:0] n6830_o;
  wire [28:0] n6831_o;
  wire [28:0] n6832_o;
  wire [28:0] n6833_o;
  wire n6835_o;
  wire [1:0] n6838_o;
  wire n6839_o;
  wire n6840_o;
  wire [4:0] n6841_o;
  wire [31:0] n6842_o;
  wire [2:0] n6843_o;
  wire [2:0] n6846_o;
  wire n6848_o;
  wire [7:0] n6849_o;
  wire [4:0] n6852_o;
  wire [2:0] n6853_o;
  wire [2:0] n6866_o;
  wire n6867_o;
  wire [1:0] n6869_o;
  wire [1:0] n6871_o;
  wire n6873_o;
  wire n6874_o;
  wire n6875_o;
  wire [3:0] n6878_o;
  wire [1:0] n6879_o;
  wire n6880_o;
  wire n6881_o;
  wire [4:0] n6883_o;
  wire [2:0] n6893_o;
  wire [2:0] n6896_o;
  wire [1:0] n6897_o;
  wire [4:0] n6898_o;
  wire n6900_o;
  wire n6901_o;
  wire n6903_o;
  wire [4:0] n6904_o;
  wire [4:0] n6905_o;
  wire [7:0] n6906_o;
  wire [7:0] n6907_o;
  wire n6909_o;
  wire n6911_o;
  wire n6912_o;
  wire [4:0] n6914_o;
  wire [2:0] n6922_o;
  wire [103:0] n6926_o;
  wire [28:0] n6927_o;
  localparam [63:0] n6933_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] n6934_o;
  wire [2:0] n6935_o;
  wire [63:0] n6936_o;
  wire [4:0] n6941_o;
  wire [2:0] n6950_o;
  wire n6951_o;
  wire [1:0] n6954_o;
  wire [1:0] n6955_o;
  wire n6956_o;
  wire n6957_o;
  wire n6958_o;
  wire [4:0] n6960_o;
  wire [2:0] n6970_o;
  wire [2:0] n6973_o;
  wire [1:0] n6974_o;
  wire [4:0] n6975_o;
  wire [4:0] n6977_o;
  wire [4:0] n6978_o;
  wire n6980_o;
  wire [2:0] n6981_o;
  reg [195:0] n6983_o;
  reg [3:0] n6985_o;
  wire [1:0] n6986_o;
  reg [1:0] n6988_o;
  wire [28:0] n6989_o;
  wire [28:0] n6990_o;
  reg [28:0] n6992_o;
  wire n6993_o;
  reg n6995_o;
  wire n6996_o;
  wire n6997_o;
  reg n6999_o;
  wire [1:0] n7000_o;
  wire [1:0] n7001_o;
  reg [1:0] n7003_o;
  wire [4:0] n7004_o;
  reg [4:0] n7006_o;
  wire [52:0] n7007_o;
  wire [48:0] n7008_o;
  wire [2:0] n7009_o;
  wire [52:0] n7010_o;
  reg [52:0] n7012_o;
  wire n7013_o;
  wire n7014_o;
  reg n7016_o;
  wire n7017_o;
  wire n7018_o;
  reg n7020_o;
  wire n7021_o;
  wire n7022_o;
  reg n7024_o;
  wire n7025_o;
  wire n7026_o;
  reg n7028_o;
  wire n7029_o;
  wire n7030_o;
  reg n7032_o;
  wire n7033_o;
  wire n7034_o;
  reg n7036_o;
  wire n7037_o;
  wire n7038_o;
  reg n7040_o;
  wire n7041_o;
  wire n7042_o;
  reg n7044_o;
  wire [195:0] n7049_o;
  wire [3:0] n7050_o;
  wire [3:0] n7051_o;
  wire [30:0] n7052_o;
  wire [1:0] n7053_o;
  wire [67:0] n7054_o;
  wire [105:0] n7055_o;
  wire [30:0] n7056_o;
  wire [30:0] n7057_o;
  wire [71:0] n7058_o;
  wire [71:0] n7059_o;
  wire [71:0] n7060_o;
  wire [1:0] n7061_o;
  wire [1:0] n7062_o;
  wire n7063_o;
  wire n7064_o;
  wire n7065_o;
  wire [67:0] n7066_o;
  wire [67:0] n7067_o;
  wire n7070_o;
  wire [1:0] n7072_o;
  wire n7074_o;
  wire n7081_o;
  wire n7082_o;
  wire n7083_o;
  wire n7085_o;
  wire n7086_o;
  wire n7087_o;
  wire n7088_o;
  wire n7089_o;
  wire n7091_o;
  wire n7092_o;
  wire n7093_o;
  wire [174:0] n7096_o;
  reg [195:0] n7115_q;
  reg [3:0] n7116_q;
  reg [3:0] n7117_q;
  wire n7118_o;
  wire n7119_o;
  wire n7120_o;
  wire n7121_o;
  wire n7124_o;
  wire n7125_o;
  wire n7126_o;
  wire n7127_o;
  reg [174:0] n7130_q;
  reg [66:0] n7131_q;
  wire [241:0] n7132_o;
  reg n7138_q;
  reg [1:0] n7139_q;
  reg n7140_q;
  wire [101:0] n7141_o;
  localparam [1:0] n7142_o = 2'bZ;
  localparam [53:0] n7143_o = 54'bZ;
  wire [63:0] n7145_data; // mem_rd
  wire [49:0] n7147_data; // mem_rd
  wire n7149_o;
  wire n7150_o;
  wire n7151_o;
  wire n7152_o;
  wire [1:0] n7153_o;
  reg n7154_o;
  wire n7155_o;
  wire n7156_o;
  wire n7157_o;
  wire n7158_o;
  wire n7159_o;
  wire n7160_o;
  wire n7161_o;
  wire n7162_o;
  wire n7163_o;
  wire n7164_o;
  wire n7165_o;
  wire n7166_o;
  wire n7167_o;
  wire n7168_o;
  wire n7169_o;
  wire n7170_o;
  wire [3:0] n7171_o;
  wire n7172_o;
  wire n7173_o;
  wire n7174_o;
  wire n7175_o;
  wire n7176_o;
  wire n7177_o;
  wire n7178_o;
  wire n7179_o;
  wire n7180_o;
  wire n7181_o;
  wire n7182_o;
  wire n7183_o;
  wire n7184_o;
  wire n7185_o;
  wire n7186_o;
  wire n7187_o;
  wire [3:0] n7188_o;
  wire n7189_o;
  wire n7190_o;
  wire n7191_o;
  wire n7192_o;
  wire [1:0] n7193_o;
  reg n7194_o;
  wire n7195_o;
  wire n7196_o;
  wire n7197_o;
  wire n7198_o;
  wire n7199_o;
  wire n7200_o;
  wire n7201_o;
  wire n7202_o;
  wire [1:0] n7203_o;
  reg n7204_o;
  wire [1:0] n7205_o;
  reg n7206_o;
  wire n7207_o;
  wire n7208_o;
  wire [48:0] n7209_o;
  wire [48:0] n7210_o;
  wire [48:0] n7211_o;
  wire [48:0] n7212_o;
  wire [1:0] n7213_o;
  reg [48:0] n7214_o;
  wire [31:0] n7215_o;
  wire [31:0] n7216_o;
  wire [31:0] n7217_o;
  wire [48:0] n7218_o;
  wire [48:0] n7219_o;
  wire [48:0] n7220_o;
  wire [48:0] n7221_o;
  wire [1:0] n7222_o;
  reg [48:0] n7223_o;
  wire n7224_o;
  wire n7225_o;
  wire n7226_o;
  wire n7227_o;
  wire n7228_o;
  wire n7229_o;
  wire n7230_o;
  wire n7231_o;
  wire n7232_o;
  wire n7233_o;
  wire n7234_o;
  wire n7235_o;
  wire n7236_o;
  wire n7237_o;
  wire n7238_o;
  wire n7239_o;
  wire [3:0] n7240_o;
  wire n7241_o;
  wire n7242_o;
  wire n7243_o;
  wire n7244_o;
  wire n7245_o;
  wire n7246_o;
  wire n7247_o;
  wire n7248_o;
  wire n7249_o;
  wire n7250_o;
  wire n7251_o;
  wire n7252_o;
  wire n7253_o;
  wire n7254_o;
  wire n7255_o;
  wire n7256_o;
  wire [3:0] n7257_o;
  wire n7258_o;
  wire n7259_o;
  wire n7260_o;
  wire n7261_o;
  wire n7262_o;
  wire n7263_o;
  wire n7264_o;
  wire n7265_o;
  wire [48:0] n7266_o;
  wire [48:0] n7267_o;
  wire [48:0] n7268_o;
  wire [48:0] n7269_o;
  wire [48:0] n7270_o;
  wire [48:0] n7271_o;
  wire [48:0] n7272_o;
  wire [48:0] n7273_o;
  wire [195:0] n7274_o;
  wire n7275_o;
  wire n7276_o;
  wire n7277_o;
  wire n7278_o;
  wire n7279_o;
  wire n7280_o;
  wire n7281_o;
  wire n7282_o;
  wire n7283_o;
  wire n7284_o;
  wire n7285_o;
  wire n7286_o;
  wire n7287_o;
  wire n7288_o;
  wire n7289_o;
  wire n7290_o;
  wire n7291_o;
  wire n7292_o;
  wire n7293_o;
  wire n7294_o;
  wire n7295_o;
  wire n7296_o;
  wire n7297_o;
  wire n7298_o;
  wire n7299_o;
  wire n7300_o;
  wire n7301_o;
  wire n7302_o;
  wire n7303_o;
  wire n7304_o;
  wire n7305_o;
  wire n7306_o;
  wire n7307_o;
  wire n7308_o;
  wire [7:0] n7309_o;
  wire n7310_o;
  wire n7311_o;
  wire n7312_o;
  wire n7313_o;
  wire n7314_o;
  wire n7315_o;
  wire n7316_o;
  wire n7317_o;
  wire n7318_o;
  wire n7319_o;
  wire n7320_o;
  wire n7321_o;
  wire n7322_o;
  wire n7323_o;
  wire n7324_o;
  wire n7325_o;
  wire [3:0] n7326_o;
  assign i_out_valid = n6289_o;
  assign i_out_stop_mark = n6290_o;
  assign i_out_fetch_failed = n6291_o;
  assign i_out_nia = n6292_o;
  assign i_out_insn = n6293_o;
  assign i_out_big_endian = n6294_o;
  assign i_out_next_predicted = n6295_o;
  assign i_out_next_pred_ntaken = n6296_o;
  assign stall_out = n6590_o;
  assign wishbone_out_adr = n6300_o;
  assign wishbone_out_dat = n6301_o;
  assign wishbone_out_sel = n6302_o;
  assign wishbone_out_cyc = n6303_o;
  assign wishbone_out_stb = n6304_o;
  assign wishbone_out_we = n6305_o;
  assign events_icache_miss = n6309_o;
  assign events_itlb_miss_resolved = n6310_o;
  assign log_out = n7143_o;
  /* fetch1.vhdl:32:9  */
  assign n6287_o = {i_in_nia, i_in_pred_ntaken, i_in_predicted, i_in_stop_mark, i_in_big_endian, i_in_priv_mode, i_in_virt_mode, i_in_req};
  assign n6289_o = n7141_o[0];
  assign n6290_o = n7141_o[1];
  /* fetch1.vhdl:153:9  */
  assign n6291_o = n7141_o[2];
  assign n6292_o = n7141_o[66:3];
  assign n6293_o = n7141_o[98:67];
  assign n6294_o = n7141_o[99];
  assign n6295_o = n7141_o[100];
  assign n6296_o = n7141_o[101];
  assign n6297_o = {m_in_pte, m_in_addr, m_in_doall, m_in_tlbie, m_in_tlbld};
  assign n6300_o = n6591_o[28:0];
  /* fetch1.vhdl:142:18  */
  assign n6301_o = n6591_o[92:29];
  assign n6302_o = n6591_o[100:93];
  assign n6303_o = n6591_o[101];
  /* fetch1.vhdl:68:18  */
  assign n6304_o = n6591_o[102];
  /* fetch1.vhdl:64:5  */
  assign n6305_o = n6591_o[103];
  /* fetch1.vhdl:66:9  */
  assign n6306_o = {wishbone_in_stall, wishbone_in_ack, wishbone_in_dat};
  assign n6307_o = {wb_snoop_in_we, wb_snoop_in_stb, wb_snoop_in_cyc, wb_snoop_in_sel, wb_snoop_in_dat, wb_snoop_in_adr};
  assign n6309_o = n7142_o[0];
  assign n6310_o = n7142_o[1];
  /* icache.vhdl:144:12  */
  assign cache_tags = n7115_q; // (signal)
  /* icache.vhdl:145:12  */
  assign cache_valids = n7116_q; // (signal)
  /* icache.vhdl:162:12  */
  assign itlb_valids = n7117_q; // (signal)
  /* icache.vhdl:169:12  */
  assign eaa_priv = n6394_o; // (signal)
  /* icache.vhdl:197:12  */
  assign r = n7132_o; // (signal)
  /* icache.vhdl:202:12  */
  assign req_index = n6480_o; // (signal)
  /* icache.vhdl:203:12  */
  assign req_row = n6488_o; // (signal)
  /* icache.vhdl:205:12  */
  assign req_tag = n6497_o; // (signal)
  /* icache.vhdl:206:12  */
  assign req_is_hit = n6550_o; // (signal)
  /* icache.vhdl:207:12  */
  assign req_is_miss = n6552_o; // (signal)
  /* icache.vhdl:208:12  */
  assign req_raddr = n6500_o; // (signal)
  /* icache.vhdl:210:12  */
  assign tlb_req_index = n6362_o; // (signal)
  /* icache.vhdl:211:12  */
  assign real_addr = n6395_o; // (signal)
  /* icache.vhdl:212:12  */
  assign ra_valid = n6397_o; // (signal)
  /* icache.vhdl:213:12  */
  assign priv_fault = n6400_o; // (signal)
  /* icache.vhdl:214:12  */
  assign access_ok = n6402_o; // (signal)
  /* icache.vhdl:558:58  */
  assign cache_out = rams_n1_dout; // (signal)
  /* icache.vhdl:226:12  */
  assign snoop_valid = n7138_q; // (signal)
  /* icache.vhdl:227:12  */
  assign snoop_index = n7139_q; // (signal)
  /* icache.vhdl:668:60  */
  assign snoop_hits = n7140_q; // (signal)
  /* icache.vhdl:365:16  */
  assign rams_n1_do_read = n6335_o; // (signal)
  /* icache.vhdl:366:16  */
  assign rams_n1_do_write = n6341_o; // (signal)
  /* icache.vhdl:367:16  */
  assign rams_n1_rd_addr = req_row; // (signal)
  /* icache.vhdl:368:16  */
  assign rams_n1_wr_addr = n6344_o; // (signal)
  /* icache.vhdl:369:16  */
  assign rams_n1_dout = rams_n1_way_rd_data; // (signal)
  /* icache.vhdl:370:16  */
  assign rams_n1_wr_sel = n6347_o; // (signal)
  /* icache.vhdl:371:16  */
  assign rams_n1_wr_dat = n6332_o; // (signal)
  /* icache.vhdl:373:9  */
  cache_ram_5_64_1489f923c4dca729178b3e3233458550d8dddf29 rams_n1_way (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(clk),
    .rd_en(rams_n1_do_read),
    .rd_addr(rams_n1_rd_addr),
    .wr_sel(rams_n1_wr_sel),
    .wr_addr(rams_n1_wr_addr),
    .wr_data(rams_n1_wr_dat),
    .rd_data(rams_n1_way_rd_data));
  /* icache.vhdl:391:27  */
  assign n6320_o = r[228];
  /* icache.vhdl:391:42  */
  assign n6321_o = ~n6320_o;
  /* icache.vhdl:392:39  */
  assign n6322_o = n6306_o[63:0];
  /* icache.vhdl:396:72  */
  assign n6323_o = n6306_o[31:24];
  /* icache.vhdl:396:72  */
  assign n6324_o = n6306_o[23:16];
  /* icache.vhdl:396:72  */
  assign n6325_o = n6306_o[15:8];
  /* icache.vhdl:396:72  */
  assign n6326_o = n6306_o[7:0];
  /* icache.vhdl:396:72  */
  assign n6327_o = n6306_o[63:56];
  /* icache.vhdl:396:72  */
  assign n6328_o = n6306_o[55:48];
  /* icache.vhdl:396:72  */
  assign n6329_o = n6306_o[47:40];
  /* icache.vhdl:396:72  */
  assign n6330_o = n6306_o[39:32];
  assign n6331_o = {n6330_o, n6329_o, n6328_o, n6327_o, n6326_o, n6325_o, n6324_o, n6323_o};
  /* icache.vhdl:391:13  */
  assign n6332_o = n6321_o ? n6322_o : n6331_o;
  /* icache.vhdl:399:24  */
  assign n6335_o = ~stall_in;
  /* icache.vhdl:401:28  */
  assign n6336_o = n6306_o[64];
  /* icache.vhdl:401:38  */
  assign n6338_o = n6336_o & 1'b1;
  /* icache.vhdl:401:13  */
  assign n6341_o = n6338_o ? 1'b1 : 1'b0;
  /* icache.vhdl:406:56  */
  assign n6344_o = r[179:175];
  assign n6347_o = {rams_n1_do_write, rams_n1_do_write, rams_n1_do_write, rams_n1_do_write, rams_n1_do_write, rams_n1_do_write, rams_n1_do_write, rams_n1_do_write};
  /* icache.vhdl:454:39  */
  assign n6352_o = n6287_o[70:7];
  /* icache.vhdl:323:21  */
  assign n6358_o = n6352_o[13:12];
  /* icache.vhdl:324:25  */
  assign n6359_o = n6352_o[15:14];
  /* icache.vhdl:324:17  */
  assign n6360_o = n6358_o ^ n6359_o;
  /* icache.vhdl:325:25  */
  assign n6361_o = n6352_o[17:16];
  /* icache.vhdl:325:17  */
  assign n6362_o = n6360_o ^ n6361_o;
  /* icache.vhdl:457:17  */
  assign n6373_o = n6287_o[1];
  /* icache.vhdl:458:29  */
  assign n6374_o = n7145_data[55:12];
  /* icache.vhdl:459:34  */
  assign n6375_o = n6287_o[18:7];
  /* icache.vhdl:458:69  */
  assign n6376_o = {n6374_o, n6375_o};
  /* icache.vhdl:460:31  */
  assign n6377_o = n6287_o[70:21];
  /* icache.vhdl:460:21  */
  assign n6378_o = n7147_data == n6377_o;
  /* icache.vhdl:461:41  */
  assign n6380_o = 2'b11 - tlb_req_index;
  /* icache.vhdl:460:13  */
  assign n6384_o = n6378_o ? n7154_o : 1'b0;
  /* icache.vhdl:465:28  */
  assign n6385_o = n7145_data[3];
  /* icache.vhdl:467:44  */
  assign n6387_o = n6287_o[70:7];
  /* common.vhdl:790:20  */
  assign n6392_o = n6387_o[55:0];
  /* icache.vhdl:457:9  */
  assign n6394_o = n6373_o ? n6385_o : 1'b1;
  /* icache.vhdl:457:9  */
  assign n6395_o = n6373_o ? n6376_o : n6392_o;
  /* icache.vhdl:457:9  */
  assign n6397_o = n6373_o ? n6384_o : 1'b1;
  /* icache.vhdl:473:45  */
  assign n6398_o = n6287_o[2];
  /* icache.vhdl:473:36  */
  assign n6399_o = ~n6398_o;
  /* icache.vhdl:473:32  */
  assign n6400_o = eaa_priv & n6399_o;
  /* icache.vhdl:474:35  */
  assign n6401_o = ~priv_fault;
  /* icache.vhdl:474:31  */
  assign n6402_o = ra_valid & n6401_o;
  /* icache.vhdl:482:38  */
  assign n6408_o = n6297_o[66:3];
  /* icache.vhdl:323:21  */
  assign n6414_o = n6408_o[13:12];
  /* icache.vhdl:324:25  */
  assign n6415_o = n6408_o[15:14];
  /* icache.vhdl:324:17  */
  assign n6416_o = n6414_o ^ n6415_o;
  /* icache.vhdl:325:25  */
  assign n6417_o = n6408_o[17:16];
  /* icache.vhdl:325:17  */
  assign n6418_o = n6416_o ^ n6417_o;
  /* icache.vhdl:483:35  */
  assign n6421_o = n6297_o[1];
  /* icache.vhdl:483:56  */
  assign n6422_o = n6297_o[2];
  /* icache.vhdl:483:47  */
  assign n6423_o = n6421_o & n6422_o;
  /* icache.vhdl:483:26  */
  assign n6424_o = rst | n6423_o;
  /* icache.vhdl:488:24  */
  assign n6429_o = n6297_o[1];
  /* icache.vhdl:490:29  */
  assign n6431_o = 2'b11 - n6418_o;
  /* icache.vhdl:491:24  */
  assign n6435_o = n6297_o[0];
  /* icache.vhdl:492:49  */
  assign n6439_o = n6297_o[66:17];
  /* icache.vhdl:493:45  */
  assign n6444_o = n6297_o[130:67];
  /* icache.vhdl:494:29  */
  assign n6447_o = 2'b11 - n6418_o;
  /* icache.vhdl:491:13  */
  assign n6451_o = n6435_o ? n7188_o : itlb_valids;
  /* icache.vhdl:488:13  */
  assign n6454_o = n6429_o ? n7171_o : n6451_o;
  assign n6457_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* icache.vhdl:483:13  */
  assign n6458_o = n6424_o ? n6457_o : n6454_o;
  /* icache.vhdl:506:37  */
  assign n6475_o = n6287_o[70:7];
  /* icache.vhdl:233:40  */
  assign n6480_o = n6475_o[7:6];
  /* icache.vhdl:507:33  */
  assign n6483_o = n6287_o[70:7];
  /* icache.vhdl:239:40  */
  assign n6488_o = n6483_o[7:3];
  /* icache.vhdl:508:44  */
  assign n6491_o = n6287_o[3];
  /* icache.vhdl:303:29  */
  assign n6496_o = real_addr[55:8];
  /* icache.vhdl:303:23  */
  assign n6497_o = {n6491_o, n6496_o};
  /* icache.vhdl:513:31  */
  assign n6498_o = real_addr[55:3];
  /* icache.vhdl:513:72  */
  assign n6500_o = {n6498_o, 3'b000};
  /* icache.vhdl:520:21  */
  assign n6501_o = n6287_o[0];
  /* icache.vhdl:521:31  */
  assign n6503_o = 2'b11 - req_index;
  /* icache.vhdl:522:21  */
  assign n6506_o = r[68:67];
  /* icache.vhdl:522:27  */
  assign n6508_o = n6506_o == 2'b11;
  /* icache.vhdl:523:29  */
  assign n6509_o = {30'b0, req_index};  //  uext
  /* icache.vhdl:523:33  */
  assign n6510_o = r[174:173];
  /* icache.vhdl:523:29  */
  assign n6511_o = {30'b0, n6510_o};  //  uext
  /* icache.vhdl:523:29  */
  assign n6512_o = n6509_o == n6511_o;
  /* icache.vhdl:522:38  */
  assign n6513_o = n6508_o & n6512_o;
  /* icache.vhdl:523:45  */
  assign n6515_o = n6513_o & 1'b1;
  /* icache.vhdl:525:40  */
  assign n6516_o = {27'b0, req_row};  //  uext
  assign n6517_o = n6516_o[2:0];
  /* icache.vhdl:525:40  */
  assign n6520_o = 3'b111 - n6517_o;
  /* icache.vhdl:524:35  */
  assign n6523_o = n6515_o & n7208_o;
  /* icache.vhdl:521:51  */
  assign n6524_o = n7194_o | n6523_o;
  /* icache.vhdl:520:31  */
  assign n6525_o = n6501_o & n6524_o;
  /* icache.vhdl:526:43  */
  assign n6528_o = 2'b11 - req_index;
  /* icache.vhdl:526:55  */
  assign n6535_o = n7214_o == req_tag;
  /* icache.vhdl:526:17  */
  assign n6538_o = n6535_o ? 1'b1 : 1'b0;
  /* icache.vhdl:520:13  */
  assign n6540_o = n6525_o ? n6538_o : 1'b0;
  /* icache.vhdl:534:17  */
  assign n6542_o = n6287_o[0];
  /* icache.vhdl:534:27  */
  assign n6543_o = n6542_o & access_ok;
  /* icache.vhdl:534:60  */
  assign n6544_o = ~flush_in;
  /* icache.vhdl:534:47  */
  assign n6545_o = n6543_o & n6544_o;
  /* icache.vhdl:534:74  */
  assign n6546_o = ~rst;
  /* icache.vhdl:534:66  */
  assign n6547_o = n6545_o & n6546_o;
  /* icache.vhdl:536:28  */
  assign n6548_o = ~n6540_o;
  /* icache.vhdl:534:9  */
  assign n6550_o = n6547_o ? n6540_o : 1'b0;
  /* icache.vhdl:534:9  */
  assign n6552_o = n6547_o ? n6548_o : 1'b0;
  /* icache.vhdl:558:40  */
  assign n6563_o = r[63:0];
  /* icache.vhdl:296:41  */
  assign n6569_o = n6563_o[2];
  /* icache.vhdl:559:26  */
  assign n6582_o = r[65];
  /* icache.vhdl:560:24  */
  assign n6583_o = r[63:0];
  /* icache.vhdl:561:30  */
  assign n6584_o = r[64];
  /* icache.vhdl:562:33  */
  assign n6585_o = r[241];
  /* icache.vhdl:563:31  */
  assign n6586_o = r[66];
  /* icache.vhdl:564:38  */
  assign n6587_o = n6287_o[5];
  /* icache.vhdl:565:40  */
  assign n6588_o = n6287_o[6];
  /* icache.vhdl:568:34  */
  assign n6589_o = n6540_o & access_ok;
  /* icache.vhdl:568:22  */
  assign n6590_o = ~n6589_o;
  /* icache.vhdl:571:27  */
  assign n6591_o = r[172:69];
  /* icache.vhdl:581:30  */
  assign n6597_o = rst | flush_in;
  assign n6599_o = r[65];
  /* icache.vhdl:581:17  */
  assign n6600_o = n6597_o ? 1'b0 : n6599_o;
  /* icache.vhdl:580:13  */
  assign n6601_o = stall_in ? n6600_o : req_is_hit;
  /* icache.vhdl:601:25  */
  assign n6602_o = ~stall_in;
  /* icache.vhdl:603:37  */
  assign n6603_o = n6287_o[4];
  /* icache.vhdl:604:35  */
  assign n6604_o = n6287_o[70:7];
  /* icache.vhdl:605:38  */
  assign n6605_o = n6287_o[3];
  assign n6606_o = {n6603_o, n6604_o};
  assign n6607_o = r[64:0];
  /* icache.vhdl:601:13  */
  assign n6608_o = n6602_o ? n6606_o : n6607_o;
  assign n6609_o = r[66];
  /* icache.vhdl:601:13  */
  assign n6610_o = n6602_o ? n6605_o : n6609_o;
  assign n6611_o = {n6610_o, n6601_o, n6608_o};
  /* icache.vhdl:643:44  */
  assign n6634_o = n6307_o[101];
  /* icache.vhdl:643:64  */
  assign n6635_o = n6307_o[102];
  /* icache.vhdl:643:48  */
  assign n6636_o = n6634_o & n6635_o;
  /* icache.vhdl:643:84  */
  assign n6637_o = n6307_o[103];
  /* icache.vhdl:643:68  */
  assign n6638_o = n6636_o & n6637_o;
  /* icache.vhdl:644:67  */
  assign n6641_o = n6307_o[28:0];
  assign n6648_o = n6647_o[63:32];
  assign n6649_o = n6647_o[2:0];
  assign n6650_o = {n6648_o, n6641_o, n6649_o};
  /* common.vhdl:790:20  */
  assign n6655_o = n6650_o[55:0];
  /* icache.vhdl:233:40  */
  assign n6661_o = n6655_o[7:6];
  /* icache.vhdl:233:40  */
  assign n6668_o = n6655_o[7:6];
  /* icache.vhdl:646:48  */
  assign n6671_o = 2'b11 - n6668_o;
  /* icache.vhdl:303:29  */
  assign n6679_o = n6655_o[55:8];
  /* icache.vhdl:303:23  */
  assign n6681_o = {1'b0, n6679_o};
  assign n6688_o = n7223_o[47:0];
  assign n6689_o = {1'b0, n6688_o};
  /* icache.vhdl:653:28  */
  assign n6690_o = n6689_o == n6681_o;
  /* icache.vhdl:653:21  */
  assign n6693_o = n6690_o ? 1'b1 : 1'b0;
  /* icache.vhdl:668:46  */
  assign n6700_o = snoop_valid & snoop_hits;
  /* icache.vhdl:669:42  */
  assign n6702_o = 2'b11 - snoop_index;
  /* icache.vhdl:668:25  */
  assign n6706_o = n6700_o ? n7240_o : cache_valids;
  assign n6707_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* icache.vhdl:659:17  */
  assign n6708_o = inval_in ? n6707_o : n6706_o;
  assign n6709_o = r[229];
  /* icache.vhdl:659:17  */
  assign n6710_o = inval_in ? 1'b0 : n6709_o;
  /* icache.vhdl:675:24  */
  assign n6711_o = r[68:67];
  /* icache.vhdl:239:40  */
  assign n6726_o = req_raddr[7:3];
  /* icache.vhdl:239:40  */
  assign n6735_o = req_raddr[7:3];
  /* icache.vhdl:247:21  */
  assign n6744_o = n6735_o[2:0];
  /* icache.vhdl:698:77  */
  assign n6746_o = n6744_o - 3'b001;
  /* wishbone_types.vhdl:69:20  */
  assign n6752_o = req_raddr[31:3];
  assign n6756_o = {n6752_o, 2'b10};
  assign n6757_o = {1'b1, 1'b1};
  assign n6758_o = {n6746_o, 1'b1, req_tag, n6726_o, req_index};
  assign n6759_o = r[97:67];
  /* icache.vhdl:683:21  */
  assign n6760_o = req_is_miss ? n6756_o : n6759_o;
  assign n6761_o = r[171:170];
  /* icache.vhdl:683:21  */
  assign n6762_o = req_is_miss ? n6757_o : n6761_o;
  assign n6763_o = r[228:173];
  assign n6764_o = r[232:230];
  assign n6765_o = {n6764_o, n6710_o, n6763_o};
  /* icache.vhdl:683:21  */
  assign n6766_o = req_is_miss ? n6758_o : n6765_o;
  /* icache.vhdl:676:17  */
  assign n6769_o = n6711_o == 2'b00;
  /* icache.vhdl:712:26  */
  assign n6770_o = r[68:67];
  /* icache.vhdl:712:32  */
  assign n6772_o = n6770_o == 2'b10;
  /* icache.vhdl:717:38  */
  assign n6774_o = 2'b11 - req_index;
  /* icache.vhdl:723:56  */
  assign n6784_o = r[228:180];
  /* icache.vhdl:724:46  */
  assign n6787_o = r[174:173];
  /* icache.vhdl:724:46  */
  assign n6789_o = 2'b11 - n6787_o;
  /* icache.vhdl:712:21  */
  assign n6793_o = n6772_o ? n7274_o : cache_tags;
  /* icache.vhdl:712:21  */
  assign n6794_o = n6772_o ? n7257_o : n6708_o;
  assign n6795_o = r[68:67];
  /* icache.vhdl:712:21  */
  assign n6796_o = n6772_o ? 2'b11 : n6795_o;
  /* icache.vhdl:732:36  */
  assign n6798_o = n6306_o[65];
  /* icache.vhdl:732:42  */
  assign n6799_o = ~n6798_o;
  /* icache.vhdl:732:54  */
  assign n6800_o = r[172:69];
  /* icache.vhdl:732:57  */
  assign n6801_o = n6800_o[102];
  /* icache.vhdl:732:48  */
  assign n6802_o = n6799_o & n6801_o;
  /* icache.vhdl:735:50  */
  assign n6804_o = r[172:69];
  /* icache.vhdl:735:53  */
  assign n6805_o = n6804_o[28:0];
  /* icache.vhdl:735:60  */
  assign n6806_o = r[232:230];
  /* icache.vhdl:253:32  */
  assign n6811_o = n6805_o[2:0];
  /* icache.vhdl:253:77  */
  assign n6812_o = n6811_o == n6806_o;
  assign n6814_o = r[171];
  /* icache.vhdl:732:21  */
  assign n6815_o = n6835_o ? 1'b0 : n6814_o;
  /* icache.vhdl:740:56  */
  assign n6817_o = r[172:69];
  /* icache.vhdl:740:59  */
  assign n6818_o = n6817_o[28:0];
  /* icache.vhdl:269:27  */
  assign n6825_o = n6818_o[2:0];
  /* icache.vhdl:270:56  */
  assign n6828_o = n6825_o + 3'b001;
  assign n6830_o = r[97:72];
  assign n6831_o = {n6830_o, n6828_o};
  assign n6832_o = r[97:69];
  /* icache.vhdl:732:21  */
  assign n6833_o = n6802_o ? n6831_o : n6832_o;
  /* icache.vhdl:732:21  */
  assign n6835_o = n6802_o & n6812_o;
  /* icache.vhdl:744:21  */
  assign n6838_o = inval_in ? 2'b01 : n6796_o;
  /* icache.vhdl:744:21  */
  assign n6839_o = inval_in ? 1'b0 : n6815_o;
  /* icache.vhdl:750:36  */
  assign n6840_o = n6306_o[64];
  /* icache.vhdl:751:40  */
  assign n6841_o = r[179:175];
  /* icache.vhdl:751:50  */
  assign n6842_o = {27'b0, n6841_o};  //  uext
  assign n6843_o = n6842_o[2:0];
  /* icache.vhdl:751:50  */
  assign n6846_o = 3'b111 - n6843_o;
  /* icache.vhdl:751:71  */
  assign n6848_o = ~inval_in;
  assign n6849_o = r[240:233];
  /* icache.vhdl:753:42  */
  assign n6852_o = r[179:175];
  /* icache.vhdl:753:55  */
  assign n6853_o = r[232:230];
  /* icache.vhdl:247:21  */
  assign n6866_o = n6852_o[2:0];
  /* icache.vhdl:259:37  */
  assign n6867_o = n6866_o == n6853_o;
  /* icache.vhdl:758:44  */
  assign n6869_o = r[174:173];
  /* icache.vhdl:758:44  */
  assign n6871_o = 2'b11 - n6869_o;
  /* icache.vhdl:758:75  */
  assign n6873_o = r[229];
  /* icache.vhdl:758:91  */
  assign n6874_o = ~inval_in;
  /* icache.vhdl:758:87  */
  assign n6875_o = n6873_o & n6874_o;
  /* icache.vhdl:750:21  */
  assign n6878_o = n6900_o ? n7326_o : n6794_o;
  /* icache.vhdl:750:21  */
  assign n6879_o = n6901_o ? 2'b00 : n6838_o;
  assign n6880_o = r[170];
  /* icache.vhdl:750:21  */
  assign n6881_o = n6903_o ? 1'b0 : n6880_o;
  /* icache.vhdl:765:51  */
  assign n6883_o = r[179:175];
  /* icache.vhdl:286:25  */
  assign n6893_o = n6883_o[2:0];
  /* icache.vhdl:287:79  */
  assign n6896_o = n6893_o + 3'b001;
  assign n6897_o = r[179:178];
  assign n6898_o = {n6897_o, n6896_o};
  /* icache.vhdl:750:21  */
  assign n6900_o = n6840_o & n6867_o;
  /* icache.vhdl:750:21  */
  assign n6901_o = n6840_o & n6867_o;
  /* icache.vhdl:750:21  */
  assign n6903_o = n6840_o & n6867_o;
  assign n6904_o = r[179:175];
  /* icache.vhdl:750:21  */
  assign n6905_o = n6840_o ? n6898_o : n6904_o;
  assign n6906_o = r[240:233];
  /* icache.vhdl:750:21  */
  assign n6907_o = n6840_o ? n7309_o : n6906_o;
  /* icache.vhdl:711:17  */
  assign n6909_o = n6711_o == 2'b10;
  /* icache.vhdl:711:30  */
  assign n6911_o = n6711_o == 2'b11;
  /* icache.vhdl:711:30  */
  assign n6912_o = n6909_o | n6911_o;
  /* icache.vhdl:771:42  */
  assign n6914_o = r[179:175];
  /* icache.vhdl:247:21  */
  assign n6922_o = n6914_o[2:0];
  /* icache.vhdl:771:92  */
  assign n6926_o = r[172:69];
  /* icache.vhdl:771:95  */
  assign n6927_o = n6926_o[28:0];
  assign n6934_o = n6933_o[63:32];
  assign n6935_o = n6933_o[2:0];
  assign n6936_o = {n6934_o, n6927_o, n6935_o};
  /* icache.vhdl:239:40  */
  assign n6941_o = n6936_o[7:3];
  /* icache.vhdl:247:21  */
  assign n6950_o = n6941_o[2:0];
  /* icache.vhdl:771:53  */
  assign n6951_o = n6922_o == n6950_o;
  assign n6954_o = r[68:67];
  /* icache.vhdl:771:21  */
  assign n6955_o = n6951_o ? 2'b00 : n6954_o;
  assign n6956_o = r[170];
  /* icache.vhdl:771:21  */
  assign n6957_o = n6951_o ? 1'b0 : n6956_o;
  /* icache.vhdl:775:36  */
  assign n6958_o = n6306_o[64];
  /* icache.vhdl:777:51  */
  assign n6960_o = r[179:175];
  /* icache.vhdl:286:25  */
  assign n6970_o = n6960_o[2:0];
  /* icache.vhdl:287:79  */
  assign n6973_o = n6970_o + 3'b001;
  assign n6974_o = r[179:178];
  assign n6975_o = {n6974_o, n6973_o};
  assign n6977_o = r[179:175];
  /* icache.vhdl:775:21  */
  assign n6978_o = n6958_o ? n6975_o : n6977_o;
  /* icache.vhdl:768:17  */
  assign n6980_o = n6711_o == 2'b01;
  assign n6981_o = {n6980_o, n6912_o, n6769_o};
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n6983_o = cache_tags;
      3'b010: n6983_o = n6793_o;
      3'b001: n6983_o = cache_tags;
      default: n6983_o = 196'bX;
    endcase
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n6985_o = n6708_o;
      3'b010: n6985_o = n6878_o;
      3'b001: n6985_o = n6708_o;
      default: n6985_o = 4'bX;
    endcase
  assign n6986_o = n6760_o[1:0];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n6988_o = n6955_o;
      3'b010: n6988_o = n6879_o;
      3'b001: n6988_o = n6986_o;
      default: n6988_o = 2'bX;
    endcase
  assign n6989_o = n6760_o[30:2];
  assign n6990_o = r[97:69];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n6992_o = n6990_o;
      3'b010: n6992_o = n6833_o;
      3'b001: n6992_o = n6989_o;
      default: n6992_o = 29'bX;
    endcase
  assign n6993_o = n6762_o[0];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n6995_o = n6957_o;
      3'b010: n6995_o = n6881_o;
      3'b001: n6995_o = n6993_o;
      default: n6995_o = 1'bX;
    endcase
  assign n6996_o = n6762_o[1];
  assign n6997_o = r[171];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n6999_o = n6997_o;
      3'b010: n6999_o = n6839_o;
      3'b001: n6999_o = n6996_o;
      default: n6999_o = 1'bX;
    endcase
  assign n7000_o = n6766_o[1:0];
  assign n7001_o = r[174:173];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n7003_o = n7001_o;
      3'b010: n7003_o = n7001_o;
      3'b001: n7003_o = n7000_o;
      default: n7003_o = 2'bX;
    endcase
  assign n7004_o = n6766_o[6:2];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n7006_o = n6978_o;
      3'b010: n7006_o = n6905_o;
      3'b001: n7006_o = n7004_o;
      default: n7006_o = 5'bX;
    endcase
  assign n7007_o = n6766_o[59:7];
  assign n7008_o = r[228:180];
  assign n7009_o = r[232:230];
  assign n7010_o = {n7009_o, n6710_o, n7008_o};
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n7012_o = n7010_o;
      3'b010: n7012_o = n7010_o;
      3'b001: n7012_o = n7007_o;
      default: n7012_o = 53'bX;
    endcase
  assign n7013_o = n6907_o[0];
  assign n7014_o = r[233];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n7016_o = n7014_o;
      3'b010: n7016_o = n7013_o;
      3'b001: n7016_o = 1'b0;
      default: n7016_o = 1'bX;
    endcase
  assign n7017_o = n6907_o[1];
  assign n7018_o = r[234];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n7020_o = n7018_o;
      3'b010: n7020_o = n7017_o;
      3'b001: n7020_o = 1'b0;
      default: n7020_o = 1'bX;
    endcase
  assign n7021_o = n6907_o[2];
  assign n7022_o = r[235];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n7024_o = n7022_o;
      3'b010: n7024_o = n7021_o;
      3'b001: n7024_o = 1'b0;
      default: n7024_o = 1'bX;
    endcase
  assign n7025_o = n6907_o[3];
  assign n7026_o = r[236];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n7028_o = n7026_o;
      3'b010: n7028_o = n7025_o;
      3'b001: n7028_o = 1'b0;
      default: n7028_o = 1'bX;
    endcase
  assign n7029_o = n6907_o[4];
  assign n7030_o = r[237];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n7032_o = n7030_o;
      3'b010: n7032_o = n7029_o;
      3'b001: n7032_o = 1'b0;
      default: n7032_o = 1'bX;
    endcase
  assign n7033_o = n6907_o[5];
  assign n7034_o = r[238];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n7036_o = n7034_o;
      3'b010: n7036_o = n7033_o;
      3'b001: n7036_o = 1'b0;
      default: n7036_o = 1'bX;
    endcase
  assign n7037_o = n6907_o[6];
  assign n7038_o = r[239];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n7040_o = n7038_o;
      3'b010: n7040_o = n7037_o;
      3'b001: n7040_o = 1'b0;
      default: n7040_o = 1'bX;
    endcase
  assign n7041_o = n6907_o[7];
  assign n7042_o = r[240];
  /* icache.vhdl:675:17  */
  always @*
    case (n6981_o)
      3'b100: n7044_o = n7042_o;
      3'b010: n7044_o = n7041_o;
      3'b001: n7044_o = 1'b0;
      default: n7044_o = 1'bX;
    endcase
  /* icache.vhdl:621:13  */
  assign n7049_o = rst ? cache_tags : n6983_o;
  assign n7050_o = {1'b0, 1'b0, 1'b0, 1'b0};
  /* icache.vhdl:621:13  */
  assign n7051_o = rst ? n7050_o : n6985_o;
  assign n7052_o = {n6992_o, n6988_o};
  assign n7053_o = {n6999_o, n6995_o};
  assign n7054_o = {n7044_o, n7040_o, n7036_o, n7032_o, n7028_o, n7024_o, n7020_o, n7016_o, n7012_o, n7006_o, n7003_o};
  assign n7055_o = {1'b0, 1'b0, 1'b0, 8'b11111111, 64'b0000000000000000000000000000000000000000000000000000000000000000, 29'b00000000000000000000000000000, 2'b00};
  assign n7056_o = n7055_o[30:0];
  /* icache.vhdl:621:13  */
  assign n7057_o = rst ? n7056_o : n7052_o;
  assign n7058_o = n7055_o[102:31];
  assign n7059_o = r[169:98];
  /* icache.vhdl:621:13  */
  assign n7060_o = rst ? n7058_o : n7059_o;
  assign n7061_o = n7055_o[104:103];
  /* icache.vhdl:621:13  */
  assign n7062_o = rst ? n7061_o : n7053_o;
  assign n7063_o = n7055_o[105];
  assign n7064_o = r[172];
  /* icache.vhdl:621:13  */
  assign n7065_o = rst ? n7063_o : n7064_o;
  assign n7066_o = r[240:173];
  /* icache.vhdl:621:13  */
  assign n7067_o = rst ? n7066_o : n7054_o;
  /* icache.vhdl:621:13  */
  assign n7070_o = rst ? 1'b0 : n6638_o;
  /* icache.vhdl:621:13  */
  assign n7072_o = rst ? 2'b00 : n6661_o;
  /* icache.vhdl:621:13  */
  assign n7074_o = rst ? 1'b0 : n6693_o;
  /* icache.vhdl:783:26  */
  assign n7081_o = rst | flush_in;
  /* icache.vhdl:783:52  */
  assign n7082_o = n6297_o[0];
  /* icache.vhdl:783:44  */
  assign n7083_o = n7081_o | n7082_o;
  /* icache.vhdl:785:24  */
  assign n7085_o = n6287_o[0];
  /* icache.vhdl:785:48  */
  assign n7086_o = ~access_ok;
  /* icache.vhdl:785:34  */
  assign n7087_o = n7085_o & n7086_o;
  /* icache.vhdl:785:67  */
  assign n7088_o = ~stall_in;
  /* icache.vhdl:785:54  */
  assign n7089_o = n7087_o & n7088_o;
  assign n7091_o = r[241];
  /* icache.vhdl:785:13  */
  assign n7092_o = n7089_o ? 1'b1 : n7091_o;
  /* icache.vhdl:783:13  */
  assign n7093_o = n7083_o ? 1'b0 : n7092_o;
  assign n7096_o = {n7093_o, n7067_o, n7065_o, n7062_o, n7060_o, n7057_o};
  /* icache.vhdl:618:9  */
  always @(posedge clk)
    n7115_q <= n7049_o;
  /* icache.vhdl:618:9  */
  always @(posedge clk)
    n7116_q <= n7051_o;
  /* icache.vhdl:481:9  */
  always @(posedge clk)
    n7117_q <= n6458_o;
  /* icache.vhdl:483:13  */
  assign n7118_o = ~n6424_o;
  /* icache.vhdl:488:13  */
  assign n7119_o = ~n6429_o;
  /* icache.vhdl:483:13  */
  assign n7120_o = n7118_o & n7119_o;
  /* icache.vhdl:483:13  */
  assign n7121_o = n7120_o & n6435_o;
  /* icache.vhdl:483:13  */
  assign n7124_o = ~n6424_o;
  /* icache.vhdl:488:13  */
  assign n7125_o = ~n6429_o;
  /* icache.vhdl:483:13  */
  assign n7126_o = n7124_o & n7125_o;
  /* icache.vhdl:483:13  */
  assign n7127_o = n7126_o & n6435_o;
  /* icache.vhdl:618:9  */
  always @(posedge clk)
    n7130_q <= n7096_o;
  /* icache.vhdl:577:9  */
  always @(posedge clk)
    n7131_q <= n6611_o;
  /* icache.vhdl:577:9  */
  assign n7132_o = {n7130_q, n7131_q};
  /* icache.vhdl:618:9  */
  always @(posedge clk)
    n7138_q <= n7070_o;
  /* icache.vhdl:618:9  */
  always @(posedge clk)
    n7139_q <= n7072_o;
  /* icache.vhdl:618:9  */
  always @(posedge clk)
    n7140_q <= n7074_o;
  /* icache.vhdl:618:9  */
  assign n7141_o = {n6588_o, n6587_o, n6586_o, n7217_o, n6583_o, n6585_o, n6584_o, n6582_o};
  /* icache.vhdl:455:26  */
  reg [63:0] itlb_ptes[3:0] ; // memory
  assign n7145_data = itlb_ptes[tlb_req_index];
  always @(posedge clk)
    if (n7127_o)
      itlb_ptes[n6418_o] <= n6444_o;
  /* icache.vhdl:455:26  */
  /* icache.vhdl:493:27  */
  /* icache.vhdl:456:27  */
  reg [49:0] itlb_tags[3:0] ; // memory
  assign n7147_data = itlb_tags[tlb_req_index];
  always @(posedge clk)
    if (n7121_o)
      itlb_tags[n6418_o] <= n6439_o;
  /* icache.vhdl:456:27  */
  /* icache.vhdl:492:27  */
  /* icache.vhdl:483:13  */
  assign n7149_o = itlb_valids[0];
  /* icache.vhdl:483:13  */
  assign n7150_o = itlb_valids[1];
  /* icache.vhdl:163:12  */
  assign n7151_o = itlb_valids[2];
  /* icache.vhdl:492:17  */
  assign n7152_o = itlb_valids[3];
  /* icache.vhdl:461:40  */
  assign n7153_o = n6380_o[1:0];
  /* icache.vhdl:461:40  */
  always @*
    case (n7153_o)
      2'b00: n7154_o = n7149_o;
      2'b01: n7154_o = n7150_o;
      2'b10: n7154_o = n7151_o;
      2'b11: n7154_o = n7152_o;
    endcase
  /* icache.vhdl:490:17  */
  assign n7155_o = n6431_o[1];
  /* icache.vhdl:490:17  */
  assign n7156_o = ~n7155_o;
  /* icache.vhdl:490:17  */
  assign n7157_o = n6431_o[0];
  /* icache.vhdl:490:17  */
  assign n7158_o = ~n7157_o;
  /* icache.vhdl:490:17  */
  assign n7159_o = n7156_o & n7158_o;
  /* icache.vhdl:490:17  */
  assign n7160_o = n7156_o & n7157_o;
  /* icache.vhdl:490:17  */
  assign n7161_o = n7155_o & n7158_o;
  /* icache.vhdl:490:17  */
  assign n7162_o = n7155_o & n7157_o;
  /* icache.vhdl:493:27  */
  assign n7163_o = itlb_valids[0];
  /* icache.vhdl:490:17  */
  assign n7164_o = n7159_o ? 1'b0 : n7163_o;
  /* icache.vhdl:382:28  */
  assign n7165_o = itlb_valids[1];
  /* icache.vhdl:490:17  */
  assign n7166_o = n7160_o ? 1'b0 : n7165_o;
  /* icache.vhdl:71:9  */
  assign n7167_o = itlb_valids[2];
  /* icache.vhdl:490:17  */
  assign n7168_o = n7161_o ? 1'b0 : n7167_o;
  /* icache.vhdl:62:9  */
  assign n7169_o = itlb_valids[3];
  /* icache.vhdl:490:17  */
  assign n7170_o = n7162_o ? 1'b0 : n7169_o;
  assign n7171_o = {n7170_o, n7168_o, n7166_o, n7164_o};
  /* icache.vhdl:494:17  */
  assign n7172_o = n6447_o[1];
  /* icache.vhdl:494:17  */
  assign n7173_o = ~n7172_o;
  /* icache.vhdl:494:17  */
  assign n7174_o = n6447_o[0];
  /* icache.vhdl:494:17  */
  assign n7175_o = ~n7174_o;
  /* icache.vhdl:494:17  */
  assign n7176_o = n7173_o & n7175_o;
  /* icache.vhdl:494:17  */
  assign n7177_o = n7173_o & n7174_o;
  /* icache.vhdl:494:17  */
  assign n7178_o = n7172_o & n7175_o;
  /* icache.vhdl:494:17  */
  assign n7179_o = n7172_o & n7174_o;
  /* icache.vhdl:618:9  */
  assign n7180_o = itlb_valids[0];
  /* icache.vhdl:494:17  */
  assign n7181_o = n7176_o ? 1'b1 : n7180_o;
  /* icache.vhdl:618:9  */
  assign n7182_o = itlb_valids[1];
  /* icache.vhdl:494:17  */
  assign n7183_o = n7177_o ? 1'b1 : n7182_o;
  assign n7184_o = itlb_valids[2];
  /* icache.vhdl:494:17  */
  assign n7185_o = n7178_o ? 1'b1 : n7184_o;
  assign n7186_o = itlb_valids[3];
  /* icache.vhdl:494:17  */
  assign n7187_o = n7179_o ? 1'b1 : n7186_o;
  /* icache.vhdl:621:13  */
  assign n7188_o = {n7187_o, n7185_o, n7183_o, n7181_o};
  /* icache.vhdl:494:29  */
  assign n7189_o = cache_valids[0];
  /* icache.vhdl:494:17  */
  assign n7190_o = cache_valids[1];
  /* icache.vhdl:621:13  */
  assign n7191_o = cache_valids[2];
  /* icache.vhdl:621:13  */
  assign n7192_o = cache_valids[3];
  /* icache.vhdl:521:41  */
  assign n7193_o = n6503_o[1:0];
  /* icache.vhdl:521:41  */
  always @*
    case (n7193_o)
      2'b00: n7194_o = n7189_o;
      2'b01: n7194_o = n7190_o;
      2'b10: n7194_o = n7191_o;
      2'b11: n7194_o = n7192_o;
    endcase
  /* icache.vhdl:521:41  */
  assign n7195_o = r[233];
  /* icache.vhdl:521:31  */
  assign n7196_o = r[234];
  /* icache.vhdl:621:13  */
  assign n7197_o = r[235];
  /* icache.vhdl:675:17  */
  assign n7198_o = r[236];
  assign n7199_o = r[237];
  /* icache.vhdl:675:17  */
  assign n7200_o = r[238];
  assign n7201_o = r[239];
  /* icache.vhdl:288:16  */
  assign n7202_o = r[240];
  /* icache.vhdl:525:31  */
  assign n7203_o = n6520_o[1:0];
  /* icache.vhdl:525:31  */
  always @*
    case (n7203_o)
      2'b00: n7204_o = n7195_o;
      2'b01: n7204_o = n7196_o;
      2'b10: n7204_o = n7197_o;
      2'b11: n7204_o = n7198_o;
    endcase
  /* icache.vhdl:525:31  */
  assign n7205_o = n6520_o[1:0];
  /* icache.vhdl:525:31  */
  always @*
    case (n7205_o)
      2'b00: n7206_o = n7199_o;
      2'b01: n7206_o = n7200_o;
      2'b10: n7206_o = n7201_o;
      2'b11: n7206_o = n7202_o;
    endcase
  /* icache.vhdl:525:31  */
  assign n7207_o = n6520_o[2];
  /* icache.vhdl:525:31  */
  assign n7208_o = n7207_o ? n7206_o : n7204_o;
  /* icache.vhdl:525:31  */
  assign n7209_o = cache_tags[48:0];
  /* icache.vhdl:525:40  */
  assign n7210_o = cache_tags[97:49];
  assign n7211_o = cache_tags[146:98];
  /* icache.vhdl:281:18  */
  assign n7212_o = cache_tags[195:147];
  /* icache.vhdl:309:22  */
  assign n7213_o = n6528_o[1:0];
  /* icache.vhdl:309:22  */
  always @*
    case (n7213_o)
      2'b00: n7214_o = n7209_o;
      2'b01: n7214_o = n7210_o;
      2'b10: n7214_o = n7211_o;
      2'b11: n7214_o = n7212_o;
    endcase
  /* icache.vhdl:309:22  */
  assign n7215_o = cache_out[31:0];
  /* icache.vhdl:526:43  */
  assign n7216_o = cache_out[63:32];
  /* icache.vhdl:297:20  */
  assign n7217_o = n6569_o ? n7216_o : n7215_o;
  /* icache.vhdl:297:20  */
  assign n7218_o = cache_tags[48:0];
  /* icache.vhdl:297:20  */
  assign n7219_o = cache_tags[97:49];
  assign n7220_o = cache_tags[146:98];
  /* icache.vhdl:280:14  */
  assign n7221_o = cache_tags[195:147];
  /* icache.vhdl:309:22  */
  assign n7222_o = n6671_o[1:0];
  /* icache.vhdl:309:22  */
  always @*
    case (n7222_o)
      2'b00: n7223_o = n7218_o;
      2'b01: n7223_o = n7219_o;
      2'b10: n7223_o = n7220_o;
      2'b11: n7223_o = n7221_o;
    endcase
  /* icache.vhdl:669:29  */
  assign n7224_o = n6702_o[1];
  /* icache.vhdl:669:29  */
  assign n7225_o = ~n7224_o;
  /* icache.vhdl:669:29  */
  assign n7226_o = n6702_o[0];
  /* icache.vhdl:669:29  */
  assign n7227_o = ~n7226_o;
  /* icache.vhdl:669:29  */
  assign n7228_o = n7225_o & n7227_o;
  /* icache.vhdl:669:29  */
  assign n7229_o = n7225_o & n7226_o;
  /* icache.vhdl:669:29  */
  assign n7230_o = n7224_o & n7227_o;
  /* icache.vhdl:669:29  */
  assign n7231_o = n7224_o & n7226_o;
  /* icache.vhdl:239:16  */
  assign n7232_o = cache_valids[0];
  /* icache.vhdl:669:29  */
  assign n7233_o = n7228_o ? 1'b0 : n7232_o;
  /* icache.vhdl:237:14  */
  assign n7234_o = cache_valids[1];
  /* icache.vhdl:669:29  */
  assign n7235_o = n7229_o ? 1'b0 : n7234_o;
  /* icache.vhdl:237:14  */
  assign n7236_o = cache_valids[2];
  /* icache.vhdl:669:29  */
  assign n7237_o = n7230_o ? 1'b0 : n7236_o;
  assign n7238_o = cache_valids[3];
  /* icache.vhdl:669:29  */
  assign n7239_o = n7231_o ? 1'b0 : n7238_o;
  /* wishbone_types.vhdl:19:14  */
  assign n7240_o = {n7239_o, n7237_o, n7235_o, n7233_o};
  /* icache.vhdl:717:25  */
  assign n7241_o = n6774_o[1];
  /* icache.vhdl:717:25  */
  assign n7242_o = ~n7241_o;
  /* icache.vhdl:717:25  */
  assign n7243_o = n6774_o[0];
  /* icache.vhdl:717:25  */
  assign n7244_o = ~n7243_o;
  /* icache.vhdl:717:25  */
  assign n7245_o = n7242_o & n7244_o;
  /* icache.vhdl:717:25  */
  assign n7246_o = n7242_o & n7243_o;
  /* icache.vhdl:717:25  */
  assign n7247_o = n7241_o & n7244_o;
  /* icache.vhdl:717:25  */
  assign n7248_o = n7241_o & n7243_o;
  /* icache.vhdl:243:14  */
  assign n7249_o = n6708_o[0];
  /* icache.vhdl:717:25  */
  assign n7250_o = n7245_o ? 1'b0 : n7249_o;
  assign n7251_o = n6708_o[1];
  /* icache.vhdl:717:25  */
  assign n7252_o = n7246_o ? 1'b0 : n7251_o;
  assign n7253_o = n6708_o[2];
  /* icache.vhdl:717:25  */
  assign n7254_o = n7247_o ? 1'b0 : n7253_o;
  assign n7255_o = n6708_o[3];
  /* icache.vhdl:717:25  */
  assign n7256_o = n7248_o ? 1'b0 : n7255_o;
  /* icache.vhdl:285:48  */
  assign n7257_o = {n7256_o, n7254_o, n7252_o, n7250_o};
  /* icache.vhdl:724:33  */
  assign n7258_o = n6789_o[1];
  /* icache.vhdl:724:33  */
  assign n7259_o = ~n7258_o;
  /* icache.vhdl:724:33  */
  assign n7260_o = n6789_o[0];
  /* icache.vhdl:724:33  */
  assign n7261_o = ~n7260_o;
  /* icache.vhdl:724:33  */
  assign n7262_o = n7259_o & n7261_o;
  /* icache.vhdl:724:33  */
  assign n7263_o = n7259_o & n7260_o;
  /* icache.vhdl:724:33  */
  assign n7264_o = n7258_o & n7261_o;
  /* icache.vhdl:724:33  */
  assign n7265_o = n7258_o & n7260_o;
  /* icache.vhdl:280:14  */
  assign n7266_o = cache_tags[48:0];
  /* icache.vhdl:724:33  */
  assign n7267_o = n7262_o ? n6784_o : n7266_o;
  assign n7268_o = cache_tags[97:49];
  /* icache.vhdl:724:33  */
  assign n7269_o = n7263_o ? n6784_o : n7268_o;
  assign n7270_o = cache_tags[146:98];
  /* icache.vhdl:724:33  */
  assign n7271_o = n7264_o ? n6784_o : n7270_o;
  /* icache.vhdl:244:18  */
  assign n7272_o = cache_tags[195:147];
  /* icache.vhdl:724:33  */
  assign n7273_o = n7265_o ? n6784_o : n7272_o;
  /* icache.vhdl:243:14  */
  assign n7274_o = {n7273_o, n7271_o, n7269_o, n7267_o};
  /* icache.vhdl:751:25  */
  assign n7275_o = n6846_o[2];
  /* icache.vhdl:751:25  */
  assign n7276_o = ~n7275_o;
  /* icache.vhdl:751:25  */
  assign n7277_o = n6846_o[1];
  /* icache.vhdl:751:25  */
  assign n7278_o = ~n7277_o;
  /* icache.vhdl:751:25  */
  assign n7279_o = n7276_o & n7278_o;
  /* icache.vhdl:751:25  */
  assign n7280_o = n7276_o & n7277_o;
  /* icache.vhdl:751:25  */
  assign n7281_o = n7275_o & n7278_o;
  /* icache.vhdl:751:25  */
  assign n7282_o = n7275_o & n7277_o;
  /* icache.vhdl:751:25  */
  assign n7283_o = n6846_o[0];
  /* icache.vhdl:751:25  */
  assign n7284_o = ~n7283_o;
  /* icache.vhdl:751:25  */
  assign n7285_o = n7279_o & n7284_o;
  /* icache.vhdl:751:25  */
  assign n7286_o = n7279_o & n7283_o;
  /* icache.vhdl:751:25  */
  assign n7287_o = n7280_o & n7284_o;
  /* icache.vhdl:751:25  */
  assign n7288_o = n7280_o & n7283_o;
  /* icache.vhdl:751:25  */
  assign n7289_o = n7281_o & n7284_o;
  /* icache.vhdl:751:25  */
  assign n7290_o = n7281_o & n7283_o;
  /* icache.vhdl:751:25  */
  assign n7291_o = n7282_o & n7284_o;
  /* icache.vhdl:751:25  */
  assign n7292_o = n7282_o & n7283_o;
  /* icache.vhdl:263:14  */
  assign n7293_o = n6849_o[0];
  /* icache.vhdl:751:25  */
  assign n7294_o = n7285_o ? n6848_o : n7293_o;
  /* icache.vhdl:263:14  */
  assign n7295_o = n6849_o[1];
  /* icache.vhdl:751:25  */
  assign n7296_o = n7286_o ? n6848_o : n7295_o;
  /* icache.vhdl:251:14  */
  assign n7297_o = n6849_o[2];
  /* icache.vhdl:751:25  */
  assign n7298_o = n7287_o ? n6848_o : n7297_o;
  /* icache.vhdl:251:14  */
  assign n7299_o = n6849_o[3];
  /* icache.vhdl:751:25  */
  assign n7300_o = n7288_o ? n6848_o : n7299_o;
  /* icache.vhdl:313:15  */
  assign n7301_o = n6849_o[4];
  /* icache.vhdl:751:25  */
  assign n7302_o = n7289_o ? n6848_o : n7301_o;
  /* icache.vhdl:722:53  */
  assign n7303_o = n6849_o[5];
  /* icache.vhdl:751:25  */
  assign n7304_o = n7290_o ? n6848_o : n7303_o;
  /* icache.vhdl:722:56  */
  assign n7305_o = n6849_o[6];
  /* icache.vhdl:751:25  */
  assign n7306_o = n7291_o ? n6848_o : n7305_o;
  /* icache.vhdl:722:56  */
  assign n7307_o = n6849_o[7];
  /* icache.vhdl:751:25  */
  assign n7308_o = n7292_o ? n6848_o : n7307_o;
  /* wishbone_types.vhdl:18:14  */
  assign n7309_o = {n7308_o, n7306_o, n7304_o, n7302_o, n7300_o, n7298_o, n7296_o, n7294_o};
  /* icache.vhdl:758:29  */
  assign n7310_o = n6871_o[1];
  /* icache.vhdl:758:29  */
  assign n7311_o = ~n7310_o;
  /* icache.vhdl:758:29  */
  assign n7312_o = n6871_o[0];
  /* icache.vhdl:758:29  */
  assign n7313_o = ~n7312_o;
  /* icache.vhdl:758:29  */
  assign n7314_o = n7311_o & n7313_o;
  /* icache.vhdl:758:29  */
  assign n7315_o = n7311_o & n7312_o;
  /* icache.vhdl:758:29  */
  assign n7316_o = n7310_o & n7313_o;
  /* icache.vhdl:758:29  */
  assign n7317_o = n7310_o & n7312_o;
  assign n7318_o = n6794_o[0];
  /* icache.vhdl:758:29  */
  assign n7319_o = n7314_o ? n6875_o : n7318_o;
  /* icache.vhdl:243:14  */
  assign n7320_o = n6794_o[1];
  /* icache.vhdl:758:29  */
  assign n7321_o = n7315_o ? n6875_o : n7320_o;
  /* icache.vhdl:243:14  */
  assign n7322_o = n6794_o[2];
  /* icache.vhdl:758:29  */
  assign n7323_o = n7316_o ? n6875_o : n7322_o;
  /* icache.vhdl:237:14  */
  assign n7324_o = n6794_o[3];
  /* icache.vhdl:758:29  */
  assign n7325_o = n7317_o ? n6875_o : n7324_o;
  assign n7326_o = {n7325_o, n7323_o, n7321_o, n7319_o};
endmodule

module fetch1_1e2926114d55612f17be0ce20b92717fa98c0d5f
  (input  clk,
   input  rst,
   input  stall_in,
   input  flush_in,
   input  inval_btc,
   input  stop_in,
   input  alt_reset_in,
   input  w_in_redirect,
   input  w_in_virt_mode,
   input  w_in_priv_mode,
   input  w_in_big_endian,
   input  w_in_mode_32bit,
   input  [63:0] w_in_redirect_nia,
   input  [63:0] w_in_br_nia,
   input  w_in_br_last,
   input  w_in_br_taken,
   input  d_in_redirect,
   input  [63:0] d_in_redirect_nia,
   output i_out_req,
   output i_out_virt_mode,
   output i_out_priv_mode,
   output i_out_big_endian,
   output i_out_stop_mark,
   output i_out_predicted,
   output i_out_pred_ntaken,
   output [63:0] i_out_nia,
   output [42:0] log_out);
  wire [134:0] n6093_o;
  wire [64:0] n6094_o;
  wire n6096_o;
  wire n6097_o;
  wire n6098_o;
  wire n6099_o;
  wire n6100_o;
  wire n6101_o;
  wire n6102_o;
  wire [63:0] n6103_o;
  wire [70:0] r;
  wire [70:0] r_next;
  wire [67:0] r_int;
  wire [67:0] r_next_int;
  wire advance_nia;
  wire [42:0] log_nia;
  reg [114:0] btc_rd_data;
  reg btc_rd_valid;
  wire n6109_o;
  wire [41:0] n6110_o;
  wire [42:0] n6111_o;
  wire n6113_o;
  wire n6114_o;
  wire n6115_o;
  wire n6116_o;
  wire n6117_o;
  wire n6118_o;
  wire n6119_o;
  wire n6120_o;
  wire n6121_o;
  wire n6122_o;
  wire [2:0] n6123_o;
  wire [2:0] n6124_o;
  wire [2:0] n6125_o;
  wire n6126_o;
  wire n6127_o;
  wire n6128_o;
  wire n6129_o;
  wire [63:0] n6130_o;
  wire n6131_o;
  wire n6132_o;
  wire [63:0] n6133_o;
  wire n6134_o;
  wire [65:0] n6135_o;
  wire [65:0] n6136_o;
  wire [65:0] n6137_o;
  wire [66:0] n6138_o;
  wire [66:0] n6139_o;
  wire [66:0] n6140_o;
  wire n6141_o;
  wire [70:0] n6142_o;
  wire [67:0] n6144_o;
  wire [4:0] n6153_o;
  wire n6162_o;
  wire [63:0] n6165_o;
  wire n6171_o;
  wire [61:0] n6172_o;
  wire [63:0] n6174_o;
  wire n6175_o;
  wire [31:0] n6177_o;
  wire [31:0] n6178_o;
  wire [31:0] n6179_o;
  wire n6180_o;
  wire n6181_o;
  wire n6182_o;
  wire n6183_o;
  wire n6184_o;
  wire [61:0] n6185_o;
  wire [63:0] n6187_o;
  wire n6188_o;
  wire [31:0] n6190_o;
  wire [31:0] n6191_o;
  wire [31:0] n6192_o;
  wire n6193_o;
  wire [63:0] n6194_o;
  wire n6197_o;
  wire [63:0] n6198_o;
  wire [63:0] n6200_o;
  wire n6201_o;
  wire [31:0] n6203_o;
  wire [31:0] n6204_o;
  wire [31:0] n6205_o;
  wire n6206_o;
  wire n6207_o;
  wire [51:0] n6208_o;
  wire [70:0] n6209_o;
  wire [51:0] n6210_o;
  wire n6211_o;
  wire n6212_o;
  wire n6213_o;
  wire n6214_o;
  wire n6215_o;
  wire [1:0] n6216_o;
  wire [1:0] n6217_o;
  wire [1:0] n6218_o;
  wire [64:0] n6219_o;
  wire n6220_o;
  wire n6221_o;
  wire n6222_o;
  wire [63:0] n6223_o;
  wire [63:0] n6224_o;
  wire [2:0] n6225_o;
  wire [2:0] n6226_o;
  wire [2:0] n6227_o;
  wire [65:0] n6228_o;
  wire [63:0] n6229_o;
  wire [1:0] n6230_o;
  wire [1:0] n6231_o;
  wire [1:0] n6232_o;
  wire [63:0] n6233_o;
  wire [63:0] n6234_o;
  wire [2:0] n6235_o;
  wire [2:0] n6236_o;
  wire [65:0] n6237_o;
  wire [2:0] n6238_o;
  wire [63:0] n6239_o;
  wire [2:0] n6240_o;
  wire [2:0] n6241_o;
  wire [1:0] n6242_o;
  wire [1:0] n6243_o;
  wire [1:0] n6244_o;
  wire [63:0] n6245_o;
  wire [63:0] n6246_o;
  wire n6247_o;
  wire [2:0] n6248_o;
  wire [2:0] n6249_o;
  wire [65:0] n6250_o;
  wire [2:0] n6251_o;
  wire [2:0] n6252_o;
  wire [1:0] n6253_o;
  wire [1:0] n6254_o;
  wire [1:0] n6255_o;
  wire [63:0] n6256_o;
  wire [63:0] n6257_o;
  wire n6258_o;
  wire n6259_o;
  wire [3:0] n6260_o;
  wire n6261_o;
  wire n6262_o;
  wire [2:0] n6263_o;
  wire [2:0] n6264_o;
  wire [2:0] n6265_o;
  wire [61:0] n6267_o;
  wire [63:0] n6269_o;
  wire n6270_o;
  wire n6271_o;
  wire n6272_o;
  wire n6273_o;
  wire n6274_o;
  wire n6275_o;
  wire n6276_o;
  wire n6277_o;
  wire n6278_o;
  wire [70:0] n6279_o;
  wire [67:0] n6280_o;
  reg [70:0] n6284_q;
  reg [67:0] n6285_q;
  reg [42:0] n6286_q;
  assign i_out_req = n6096_o;
  assign i_out_virt_mode = n6097_o;
  assign i_out_priv_mode = n6098_o;
  assign i_out_big_endian = n6099_o;
  assign i_out_stop_mark = n6100_o;
  assign i_out_predicted = n6101_o;
  assign i_out_pred_ntaken = n6102_o;
  assign i_out_nia = n6103_o;
  assign log_out = log_nia;
  /* wishbone_debug_master.vhdl:18:10  */
  assign n6093_o = {w_in_br_taken, w_in_br_last, w_in_br_nia, w_in_redirect_nia, w_in_mode_32bit, w_in_big_endian, w_in_priv_mode, w_in_virt_mode, w_in_redirect};
  /* wishbone_debug_master.vhdl:15:10  */
  assign n6094_o = {d_in_redirect_nia, d_in_redirect};
  assign n6096_o = r[0];
  /* wishbone_debug_master.vhdl:143:5  */
  assign n6097_o = r[1];
  assign n6098_o = r[2];
  /* wishbone_debug_master.vhdl:135:9  */
  assign n6099_o = r[3];
  /* wishbone_debug_master.vhdl:133:5  */
  assign n6100_o = r[4];
  assign n6101_o = r[5];
  /* wishbone_debug_master.vhdl:70:18  */
  assign n6102_o = r[6];
  /* wishbone_debug_master.vhdl:70:18  */
  assign n6103_o = r[70:7];
  /* fetch1.vhdl:47:12  */
  assign r = n6284_q; // (signal)
  /* fetch1.vhdl:47:15  */
  assign r_next = n6279_o; // (signal)
  /* fetch1.vhdl:48:12  */
  assign r_int = n6285_q; // (signal)
  /* fetch1.vhdl:48:19  */
  assign r_next_int = n6280_o; // (signal)
  /* fetch1.vhdl:49:12  */
  assign advance_nia = n6278_o; // (signal)
  /* fetch1.vhdl:50:12  */
  assign log_nia = n6286_q; // (signal)
  /* fetch1.vhdl:59:12  */
  always @*
    btc_rd_data = 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // (isignal)
  initial
    btc_rd_data = 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* fetch1.vhdl:60:12  */
  always @*
    btc_rd_valid = 1'b0; // (isignal)
  initial
    btc_rd_valid = 1'b0;
  /* fetch1.vhdl:67:29  */
  assign n6109_o = r[70];
  /* fetch1.vhdl:67:41  */
  assign n6110_o = r[50:9];
  /* fetch1.vhdl:67:34  */
  assign n6111_o = {n6109_o, n6110_o};
  /* fetch1.vhdl:79:34  */
  assign n6113_o = n6093_o[0];
  /* fetch1.vhdl:79:26  */
  assign n6114_o = rst | n6113_o;
  /* fetch1.vhdl:79:57  */
  assign n6115_o = n6094_o[0];
  /* fetch1.vhdl:79:49  */
  assign n6116_o = n6114_o | n6115_o;
  /* fetch1.vhdl:79:84  */
  assign n6117_o = ~stall_in;
  /* fetch1.vhdl:79:72  */
  assign n6118_o = n6116_o | n6117_o;
  /* fetch1.vhdl:80:39  */
  assign n6119_o = r_next[1];
  /* fetch1.vhdl:81:39  */
  assign n6120_o = r_next[2];
  /* fetch1.vhdl:82:40  */
  assign n6121_o = r_next[3];
  /* fetch1.vhdl:83:48  */
  assign n6122_o = r_next_int[0];
  assign n6123_o = {n6121_o, n6120_o, n6119_o};
  assign n6124_o = r[3:1];
  /* fetch1.vhdl:79:13  */
  assign n6125_o = n6118_o ? n6123_o : n6124_o;
  assign n6126_o = r_int[0];
  /* fetch1.vhdl:79:13  */
  assign n6127_o = n6118_o ? n6122_o : n6126_o;
  /* fetch1.vhdl:86:39  */
  assign n6128_o = r_next[5];
  /* fetch1.vhdl:87:41  */
  assign n6129_o = r_next[6];
  /* fetch1.vhdl:88:33  */
  assign n6130_o = r_next[70:7];
  /* fetch1.vhdl:89:53  */
  assign n6131_o = r_next_int[2];
  /* fetch1.vhdl:90:52  */
  assign n6132_o = r_next_int[3];
  /* fetch1.vhdl:91:51  */
  assign n6133_o = r_next_int[67:4];
  /* fetch1.vhdl:92:49  */
  assign n6134_o = r_next_int[1];
  assign n6135_o = {n6130_o, n6129_o, n6128_o};
  assign n6136_o = r[70:5];
  /* fetch1.vhdl:85:13  */
  assign n6137_o = advance_nia ? n6135_o : n6136_o;
  assign n6138_o = {n6133_o, n6132_o, n6131_o, n6134_o};
  assign n6139_o = r_int[67:1];
  /* fetch1.vhdl:85:13  */
  assign n6140_o = advance_nia ? n6138_o : n6139_o;
  /* fetch1.vhdl:96:22  */
  assign n6141_o = ~rst;
  assign n6142_o = {n6137_o, stop_in, n6125_o, n6141_o};
  assign n6144_o = {n6140_o, n6127_o};
  assign n6153_o = r[4:0];
  assign n6162_o = r_int[0];
  /* fetch1.vhdl:154:13  */
  assign n6165_o = alt_reset_in ? 64'b1111111111111111111111111111111111110000000000000000000000000000 : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* fetch1.vhdl:164:20  */
  assign n6171_o = n6093_o[0];
  /* fetch1.vhdl:165:39  */
  assign n6172_o = n6093_o[68:7];
  /* fetch1.vhdl:165:53  */
  assign n6174_o = {n6172_o, 2'b00};
  /* fetch1.vhdl:166:21  */
  assign n6175_o = n6093_o[4];
  assign n6177_o = n6174_o[63:32];
  /* fetch1.vhdl:166:13  */
  assign n6178_o = n6175_o ? 32'b00000000000000000000000000000000 : n6177_o;
  assign n6179_o = n6174_o[31:0];
  /* fetch1.vhdl:169:33  */
  assign n6180_o = n6093_o[1];
  /* fetch1.vhdl:170:33  */
  assign n6181_o = n6093_o[2];
  /* fetch1.vhdl:171:34  */
  assign n6182_o = n6093_o[3];
  /* fetch1.vhdl:172:38  */
  assign n6183_o = n6093_o[4];
  /* fetch1.vhdl:173:20  */
  assign n6184_o = n6094_o[0];
  /* fetch1.vhdl:174:39  */
  assign n6185_o = n6094_o[64:3];
  /* fetch1.vhdl:174:53  */
  assign n6187_o = {n6185_o, 2'b00};
  /* fetch1.vhdl:175:22  */
  assign n6188_o = r_int[0];
  assign n6190_o = n6187_o[63:32];
  /* fetch1.vhdl:175:13  */
  assign n6191_o = n6188_o ? 32'b00000000000000000000000000000000 : n6190_o;
  assign n6192_o = n6187_o[31:0];
  /* fetch1.vhdl:178:21  */
  assign n6193_o = r_int[2];
  /* fetch1.vhdl:179:28  */
  assign n6194_o = r_int[67:4];
  /* fetch1.vhdl:183:36  */
  assign n6197_o = r_int[3];
  /* fetch1.vhdl:184:51  */
  assign n6198_o = r[70:7];
  /* fetch1.vhdl:184:56  */
  assign n6200_o = n6198_o + 64'b0000000000000000000000000000000000000000000000000000000000000100;
  /* fetch1.vhdl:185:22  */
  assign n6201_o = r_int[0];
  assign n6203_o = n6200_o[63:32];
  /* fetch1.vhdl:185:13  */
  assign n6204_o = n6201_o ? 32'b00000000000000000000000000000000 : n6203_o;
  assign n6205_o = n6200_o[31:0];
  /* fetch1.vhdl:188:45  */
  assign n6206_o = r_int[1];
  /* fetch1.vhdl:188:35  */
  assign n6207_o = btc_rd_valid & n6206_o;
  /* fetch1.vhdl:189:28  */
  assign n6208_o = btc_rd_data[113:62];
  assign n6209_o = {n6204_o, n6205_o, n6197_o, 1'b0, n6153_o};
  /* fetch1.vhdl:190:24  */
  assign n6210_o = n6209_o[70:19];
  /* fetch1.vhdl:190:17  */
  assign n6211_o = n6208_o == n6210_o;
  /* fetch1.vhdl:188:63  */
  assign n6212_o = n6207_o & n6211_o;
  /* fetch1.vhdl:191:53  */
  assign n6213_o = btc_rd_data[114];
  /* fetch1.vhdl:192:56  */
  assign n6214_o = btc_rd_data[114];
  /* fetch1.vhdl:192:41  */
  assign n6215_o = ~n6214_o;
  assign n6216_o = {n6215_o, n6213_o};
  assign n6217_o = {1'b0, 1'b0};
  /* fetch1.vhdl:188:13  */
  assign n6218_o = n6212_o ? n6216_o : n6217_o;
  assign n6219_o = {n6204_o, n6205_o, n6197_o};
  /* fetch1.vhdl:178:9  */
  assign n6220_o = n6193_o ? 1'b1 : 1'b0;
  assign n6221_o = n6219_o[0];
  /* fetch1.vhdl:178:9  */
  assign n6222_o = n6193_o ? 1'b0 : n6221_o;
  assign n6223_o = n6219_o[64:1];
  /* fetch1.vhdl:178:9  */
  assign n6224_o = n6193_o ? n6194_o : n6223_o;
  assign n6225_o = {n6218_o, 1'b1};
  assign n6226_o = {1'b0, 1'b0, 1'b0};
  /* fetch1.vhdl:178:9  */
  assign n6227_o = n6193_o ? n6226_o : n6225_o;
  assign n6228_o = {n6224_o, n6222_o, n6220_o};
  assign n6229_o = {n6191_o, n6192_o};
  assign n6230_o = n6228_o[1:0];
  assign n6231_o = {1'b0, 1'b0};
  /* fetch1.vhdl:173:9  */
  assign n6232_o = n6184_o ? n6231_o : n6230_o;
  assign n6233_o = n6228_o[65:2];
  /* fetch1.vhdl:173:9  */
  assign n6234_o = n6184_o ? n6229_o : n6233_o;
  assign n6235_o = {1'b0, 1'b0, 1'b0};
  /* fetch1.vhdl:173:9  */
  assign n6236_o = n6184_o ? n6235_o : n6227_o;
  assign n6237_o = {n6234_o, n6232_o};
  assign n6238_o = {n6182_o, n6181_o, n6180_o};
  assign n6239_o = {n6178_o, n6179_o};
  assign n6240_o = r[3:1];
  /* fetch1.vhdl:164:9  */
  assign n6241_o = n6171_o ? n6238_o : n6240_o;
  assign n6242_o = n6237_o[1:0];
  assign n6243_o = {1'b0, 1'b0};
  /* fetch1.vhdl:164:9  */
  assign n6244_o = n6171_o ? n6243_o : n6242_o;
  assign n6245_o = n6237_o[65:2];
  /* fetch1.vhdl:164:9  */
  assign n6246_o = n6171_o ? n6239_o : n6245_o;
  /* fetch1.vhdl:164:9  */
  assign n6247_o = n6171_o ? n6183_o : n6162_o;
  assign n6248_o = {1'b0, 1'b0, 1'b0};
  /* fetch1.vhdl:164:9  */
  assign n6249_o = n6171_o ? n6248_o : n6236_o;
  assign n6250_o = {n6246_o, n6244_o};
  assign n6251_o = {1'b0, 1'b1, 1'b0};
  /* fetch1.vhdl:153:9  */
  assign n6252_o = rst ? n6251_o : n6241_o;
  assign n6253_o = n6250_o[1:0];
  assign n6254_o = {1'b0, 1'b0};
  /* fetch1.vhdl:153:9  */
  assign n6255_o = rst ? n6254_o : n6253_o;
  assign n6256_o = n6250_o[65:2];
  /* fetch1.vhdl:153:9  */
  assign n6257_o = rst ? n6165_o : n6256_o;
  assign n6258_o = r[4];
  assign n6259_o = r[0];
  assign n6260_o = {n6249_o, n6247_o};
  assign n6261_o = n6260_o[0];
  /* fetch1.vhdl:153:9  */
  assign n6262_o = rst ? 1'b0 : n6261_o;
  assign n6263_o = n6260_o[3:1];
  assign n6264_o = {1'b0, 1'b0, 1'b0};
  /* fetch1.vhdl:153:9  */
  assign n6265_o = rst ? n6264_o : n6263_o;
  /* fetch1.vhdl:195:43  */
  assign n6267_o = btc_rd_data[61:0];
  /* fetch1.vhdl:195:74  */
  assign n6269_o = {n6267_o, 2'b00};
  /* fetch1.vhdl:199:36  */
  assign n6270_o = n6093_o[0];
  /* fetch1.vhdl:199:28  */
  assign n6271_o = rst | n6270_o;
  /* fetch1.vhdl:199:53  */
  assign n6272_o = n6094_o[0];
  /* fetch1.vhdl:199:45  */
  assign n6273_o = n6271_o | n6272_o;
  /* fetch1.vhdl:199:72  */
  assign n6274_o = r[4];
  /* fetch1.vhdl:199:66  */
  assign n6275_o = ~n6274_o;
  /* fetch1.vhdl:199:86  */
  assign n6276_o = ~stall_in;
  /* fetch1.vhdl:199:82  */
  assign n6277_o = n6275_o & n6276_o;
  /* fetch1.vhdl:199:62  */
  assign n6278_o = n6273_o | n6277_o;
  assign n6279_o = {n6257_o, n6255_o, n6258_o, n6252_o, n6259_o};
  assign n6280_o = {n6269_o, n6265_o, n6262_o};
  /* fetch1.vhdl:66:9  */
  always @(posedge clk)
    n6284_q <= n6142_o;
  /* fetch1.vhdl:66:9  */
  always @(posedge clk)
    n6285_q <= n6144_o;
  /* fetch1.vhdl:66:9  */
  always @(posedge clk)
    n6286_q <= n6111_o;
endmodule

module wishbone_debug_master
  (input  clk,
   input  rst,
   input  [1:0] dmi_addr,
   input  [63:0] dmi_din,
   input  dmi_req,
   input  dmi_wr,
   input  [63:0] wb_in_dat,
   input  wb_in_ack,
   input  wb_in_stall,
   output [63:0] dmi_dout,
   output dmi_ack,
   output [28:0] wb_out_adr,
   output [63:0] wb_out_dat,
   output [7:0] wb_out_sel,
   output wb_out_cyc,
   output wb_out_stb,
   output wb_out_we);
  wire [28:0] n5874_o;
  wire [63:0] n5875_o;
  wire [7:0] n5876_o;
  wire n5877_o;
  wire n5878_o;
  wire n5879_o;
  wire [65:0] n5880_o;
  wire [63:0] reg_addr;
  wire [63:0] reg_ctrl_out;
  wire [10:0] reg_ctrl;
  wire [63:0] data_latch;
  wire [1:0] state;
  wire do_inc;
  wire [3:0] n5934_o;
  wire [3:0] n5935_o;
  wire [3:0] n5936_o;
  wire [3:0] n5937_o;
  wire [3:0] n5938_o;
  wire [3:0] n5939_o;
  wire [3:0] n5940_o;
  wire [3:0] n5941_o;
  wire [3:0] n5942_o;
  wire [3:0] n5943_o;
  wire [3:0] n5944_o;
  wire [3:0] n5945_o;
  wire [3:0] n5946_o;
  wire [11:0] n5947_o;
  wire [15:0] n5948_o;
  wire [15:0] n5949_o;
  wire [15:0] n5950_o;
  wire [15:0] n5951_o;
  wire [63:0] n5952_o;
  wire n5954_o;
  wire n5956_o;
  wire n5958_o;
  wire [2:0] n5960_o;
  reg [63:0] n5961_o;
  wire [1:0] n5965_o;
  wire n5972_o;
  wire n5975_o;
  wire n5978_o;
  wire n5981_o;
  wire [3:0] n5983_o;
  reg [3:0] n5984_o;
  wire [30:0] n5985_o;
  wire [63:0] n5986_o;
  wire [63:0] n5987_o;
  wire n5988_o;
  wire n5990_o;
  wire n5992_o;
  wire [10:0] n5993_o;
  wire [10:0] n5994_o;
  wire [63:0] n5995_o;
  wire [10:0] n5996_o;
  wire n5997_o;
  wire [10:0] n5998_o;
  wire [63:0] n5999_o;
  wire [10:0] n6000_o;
  wire [63:0] n6002_o;
  wire [10:0] n6004_o;
  wire n6009_o;
  wire n6011_o;
  wire n6012_o;
  wire n6013_o;
  wire [28:0] n6015_o;
  wire [7:0] n6016_o;
  wire n6019_o;
  wire n6020_o;
  wire n6025_o;
  wire n6026_o;
  wire n6027_o;
  wire n6028_o;
  wire n6029_o;
  wire [63:0] n6030_o;
  wire n6038_o;
  wire n6039_o;
  wire n6041_o;
  wire n6042_o;
  wire [1:0] n6044_o;
  wire n6046_o;
  wire n6047_o;
  wire n6048_o;
  wire n6050_o;
  wire n6051_o;
  wire n6052_o;
  wire n6054_o;
  wire n6055_o;
  wire [1:0] n6057_o;
  wire n6058_o;
  wire n6060_o;
  wire n6061_o;
  wire [1:0] n6063_o;
  wire n6065_o;
  wire [2:0] n6066_o;
  wire n6067_o;
  reg n6069_o;
  reg [1:0] n6071_o;
  reg n6074_o;
  wire n6075_o;
  wire [1:0] n6077_o;
  wire n6079_o;
  reg [63:0] n6085_q;
  reg [10:0] n6086_q;
  wire [63:0] n6087_o;
  reg [63:0] n6088_q;
  reg [1:0] n6089_q;
  reg n6090_q;
  reg n6091_q;
  wire [103:0] n6092_o;
  assign dmi_dout = n5961_o;
  assign dmi_ack = n6013_o;
  assign wb_out_adr = n5874_o;
  assign wb_out_dat = n5875_o;
  assign wb_out_sel = n5876_o;
  assign wb_out_cyc = n5877_o;
  assign wb_out_stb = n5878_o;
  assign wb_out_we = n5879_o;
  /* dmi_dtm_jtag.vhdl:175:40  */
  assign n5874_o = n6092_o[28:0];
  /* dmi_dtm_jtag.vhdl:172:40  */
  assign n5875_o = n6092_o[92:29];
  /* dmi_dtm_jtag.vhdl:81:10  */
  assign n5876_o = n6092_o[100:93];
  /* dmi_dtm_jtag.vhdl:74:10  */
  assign n5877_o = n6092_o[101];
  /* dmi_dtm_jtag.vhdl:73:10  */
  assign n5878_o = n6092_o[102];
  /* dmi_dtm_jtag.vhdl:72:10  */
  assign n5879_o = n6092_o[103];
  /* dmi_dtm_jtag.vhdl:70:10  */
  assign n5880_o = {wb_in_stall, wb_in_ack, wb_in_dat};
  /* wishbone_debug_master.vhdl:45:12  */
  assign reg_addr = n6085_q; // (signal)
  /* wishbone_debug_master.vhdl:46:12  */
  assign reg_ctrl_out = n5952_o; // (signal)
  /* wishbone_debug_master.vhdl:47:12  */
  assign reg_ctrl = n6086_q; // (signal)
  /* wishbone_debug_master.vhdl:48:12  */
  assign data_latch = n6088_q; // (signal)
  /* wishbone_debug_master.vhdl:51:12  */
  assign state = n6089_q; // (signal)
  /* wishbone_debug_master.vhdl:52:12  */
  assign do_inc = n6090_q; // (signal)
  assign n5934_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5935_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5936_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5937_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5938_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5939_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5940_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5941_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5942_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5943_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5944_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5945_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5946_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n5947_o = {1'b0, reg_ctrl};
  assign n5948_o = {n5934_o, n5935_o, n5936_o, n5937_o};
  assign n5949_o = {n5938_o, n5939_o, n5940_o, n5941_o};
  assign n5950_o = {n5942_o, n5943_o, n5944_o, n5945_o};
  assign n5951_o = {n5946_o, n5947_o};
  assign n5952_o = {n5948_o, n5949_o, n5950_o, n5951_o};
  /* wishbone_debug_master.vhdl:62:25  */
  assign n5954_o = dmi_addr == 2'b00;
  /* wishbone_debug_master.vhdl:63:25  */
  assign n5956_o = dmi_addr == 2'b01;
  /* wishbone_debug_master.vhdl:64:25  */
  assign n5958_o = dmi_addr == 2'b10;
  assign n5960_o = {n5958_o, n5956_o, n5954_o};
  /* wishbone_debug_master.vhdl:61:5  */
  always @*
    case (n5960_o)
      3'b100: n5961_o = reg_ctrl_out;
      3'b010: n5961_o = data_latch;
      3'b001: n5961_o = reg_addr;
      default: n5961_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* wishbone_debug_master.vhdl:91:74  */
  assign n5965_o = reg_ctrl[10:9];
  /* wishbone_debug_master.vhdl:74:13  */
  assign n5972_o = n5965_o == 2'b00;
  /* wishbone_debug_master.vhdl:75:13  */
  assign n5975_o = n5965_o == 2'b01;
  /* wishbone_debug_master.vhdl:76:13  */
  assign n5978_o = n5965_o == 2'b10;
  /* wishbone_debug_master.vhdl:77:13  */
  assign n5981_o = n5965_o == 2'b11;
  assign n5983_o = {n5981_o, n5978_o, n5975_o, n5972_o};
  /* wishbone_debug_master.vhdl:73:13  */
  always @*
    case (n5983_o)
      4'b1000: n5984_o = 4'b1000;
      4'b0100: n5984_o = 4'b0100;
      4'b0010: n5984_o = 4'b0010;
      4'b0001: n5984_o = 4'b0001;
      default: n5984_o = 4'b1000;
    endcase
  /* wishbone_debug_master.vhdl:90:70  */
  assign n5985_o = {27'b0, n5984_o};  //  uext
  /* wishbone_debug_master.vhdl:90:70  */
  assign n5986_o = {33'b0, n5985_o};  //  uext
  /* wishbone_debug_master.vhdl:90:70  */
  assign n5987_o = reg_addr + n5986_o;
  /* wishbone_debug_master.vhdl:92:31  */
  assign n5988_o = dmi_req & dmi_wr;
  /* wishbone_debug_master.vhdl:93:33  */
  assign n5990_o = dmi_addr == 2'b00;
  /* wishbone_debug_master.vhdl:95:36  */
  assign n5992_o = dmi_addr == 2'b10;
  /* wishbone_debug_master.vhdl:96:44  */
  assign n5993_o = dmi_din[10:0];
  /* wishbone_debug_master.vhdl:95:21  */
  assign n5994_o = n5992_o ? n5993_o : reg_ctrl;
  /* wishbone_debug_master.vhdl:92:17  */
  assign n5995_o = n5997_o ? dmi_din : reg_addr;
  /* wishbone_debug_master.vhdl:93:21  */
  assign n5996_o = n5990_o ? reg_ctrl : n5994_o;
  /* wishbone_debug_master.vhdl:92:17  */
  assign n5997_o = n5988_o & n5990_o;
  /* wishbone_debug_master.vhdl:92:17  */
  assign n5998_o = n5988_o ? n5996_o : reg_ctrl;
  /* wishbone_debug_master.vhdl:88:17  */
  assign n5999_o = do_inc ? n5987_o : n5995_o;
  /* wishbone_debug_master.vhdl:88:17  */
  assign n6000_o = do_inc ? reg_ctrl : n5998_o;
  /* wishbone_debug_master.vhdl:84:13  */
  assign n6002_o = rst ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : n5999_o;
  /* wishbone_debug_master.vhdl:84:13  */
  assign n6004_o = rst ? 11'b00000000000 : n6000_o;
  /* wishbone_debug_master.vhdl:118:39  */
  assign n6009_o = dmi_addr != 2'b01;
  /* wishbone_debug_master.vhdl:118:63  */
  assign n6011_o = state == 2'b10;
  /* wishbone_debug_master.vhdl:118:54  */
  assign n6012_o = n6009_o | n6011_o;
  /* wishbone_debug_master.vhdl:118:24  */
  assign n6013_o = n6012_o ? dmi_req : 1'b0;
  /* wishbone_debug_master.vhdl:121:27  */
  assign n6015_o = reg_addr[31:3];
  /* wishbone_debug_master.vhdl:123:27  */
  assign n6016_o = reg_ctrl[7:0];
  /* wishbone_debug_master.vhdl:127:34  */
  assign n6019_o = state == 2'b01;
  /* wishbone_debug_master.vhdl:127:23  */
  assign n6020_o = n6019_o ? 1'b1 : 1'b0;
  /* wishbone_debug_master.vhdl:136:22  */
  assign n6025_o = state == 2'b01;
  /* wishbone_debug_master.vhdl:136:43  */
  assign n6026_o = n5880_o[64];
  /* wishbone_debug_master.vhdl:136:33  */
  assign n6027_o = n6025_o & n6026_o;
  /* wishbone_debug_master.vhdl:136:64  */
  assign n6028_o = ~dmi_wr;
  /* wishbone_debug_master.vhdl:136:53  */
  assign n6029_o = n6027_o & n6028_o;
  /* wishbone_debug_master.vhdl:137:37  */
  assign n6030_o = n5880_o[63:0];
  /* wishbone_debug_master.vhdl:153:51  */
  assign n6038_o = dmi_addr == 2'b01;
  /* wishbone_debug_master.vhdl:153:38  */
  assign n6039_o = dmi_req & n6038_o;
  assign n6041_o = n6092_o[102];
  /* wishbone_debug_master.vhdl:153:21  */
  assign n6042_o = n6039_o ? 1'b1 : n6041_o;
  /* wishbone_debug_master.vhdl:153:21  */
  assign n6044_o = n6039_o ? 2'b01 : state;
  /* wishbone_debug_master.vhdl:152:17  */
  assign n6046_o = state == 2'b00;
  /* wishbone_debug_master.vhdl:158:30  */
  assign n6047_o = n5880_o[65];
  /* wishbone_debug_master.vhdl:158:36  */
  assign n6048_o = ~n6047_o;
  assign n6050_o = n6092_o[102];
  /* wishbone_debug_master.vhdl:158:21  */
  assign n6051_o = n6048_o ? 1'b0 : n6050_o;
  /* wishbone_debug_master.vhdl:161:30  */
  assign n6052_o = n5880_o[64];
  /* wishbone_debug_master.vhdl:167:43  */
  assign n6054_o = reg_ctrl[8];
  /* wishbone_debug_master.vhdl:161:21  */
  assign n6055_o = n6052_o ? 1'b0 : n6051_o;
  /* wishbone_debug_master.vhdl:161:21  */
  assign n6057_o = n6052_o ? 2'b10 : state;
  /* wishbone_debug_master.vhdl:161:21  */
  assign n6058_o = n6052_o ? n6054_o : do_inc;
  /* wishbone_debug_master.vhdl:157:17  */
  assign n6060_o = state == 2'b01;
  /* wishbone_debug_master.vhdl:170:32  */
  assign n6061_o = ~dmi_req;
  /* wishbone_debug_master.vhdl:170:21  */
  assign n6063_o = n6061_o ? 2'b00 : state;
  /* wishbone_debug_master.vhdl:169:17  */
  assign n6065_o = state == 2'b10;
  assign n6066_o = {n6065_o, n6060_o, n6046_o};
  assign n6067_o = n6092_o[102];
  /* wishbone_debug_master.vhdl:151:17  */
  always @*
    case (n6066_o)
      3'b100: n6069_o = n6067_o;
      3'b010: n6069_o = n6055_o;
      3'b001: n6069_o = n6042_o;
      default: n6069_o = 1'bX;
    endcase
  /* wishbone_debug_master.vhdl:151:17  */
  always @*
    case (n6066_o)
      3'b100: n6071_o = n6063_o;
      3'b010: n6071_o = n6057_o;
      3'b001: n6071_o = n6044_o;
      default: n6071_o = 2'bX;
    endcase
  /* wishbone_debug_master.vhdl:151:17  */
  always @*
    case (n6066_o)
      3'b100: n6074_o = 1'b0;
      3'b010: n6074_o = n6058_o;
      3'b001: n6074_o = do_inc;
      default: n6074_o = 1'bX;
    endcase
  /* wishbone_debug_master.vhdl:146:13  */
  assign n6075_o = rst ? 1'b0 : n6069_o;
  /* wishbone_debug_master.vhdl:146:13  */
  assign n6077_o = rst ? 2'b00 : n6071_o;
  /* wishbone_debug_master.vhdl:146:13  */
  assign n6079_o = rst ? 1'b0 : n6074_o;
  /* wishbone_debug_master.vhdl:83:9  */
  always @(posedge clk)
    n6085_q <= n6002_o;
  /* wishbone_debug_master.vhdl:83:9  */
  always @(posedge clk)
    n6086_q <= n6004_o;
  /* wishbone_debug_master.vhdl:135:9  */
  assign n6087_o = n6029_o ? n6030_o : data_latch;
  /* wishbone_debug_master.vhdl:135:9  */
  always @(posedge clk)
    n6088_q <= n6087_o;
  /* wishbone_debug_master.vhdl:145:9  */
  always @(posedge clk)
    n6089_q <= n6077_o;
  /* wishbone_debug_master.vhdl:145:9  */
  always @(posedge clk)
    n6090_q <= n6079_o;
  /* wishbone_debug_master.vhdl:145:9  */
  always @(posedge clk)
    n6091_q <= n6075_o;
  /* wishbone_debug_master.vhdl:145:9  */
  assign n6092_o = {dmi_wr, n6091_q, n6020_o, n6016_o, dmi_din, n6015_o};
endmodule

module dmi_dtm_jtag_8_64
  (input  sys_clk,
   input  sys_reset,
   input  [63:0] dmi_din,
   input  dmi_ack,
   input  jtag_tck,
   input  jtag_tdi,
   input  jtag_tms,
   input  jtag_trst,
   output [7:0] dmi_addr,
   output [63:0] dmi_dout,
   output dmi_req,
   output dmi_wr,
   output jtag_tdo);
  wire capture;
  wire update;
  wire sel;
  wire shift;
  wire tdi;
  wire tdo;
  wire [73:0] shiftr;
  wire [73:0] request;
  wire jtag_req;
  wire dmi_ack_0;
  wire dmi_ack_1;
  wire jtag_req_0;
  wire jtag_req_1;
  wire jtag_bsy;
  wire op_valid;
  wire [1:0] rsp_op;
  wire tap_top0_tdo_pad_o;
  wire tap_top0_tdo_padoe_o;
  wire tap_top0_shift_dr_o;
  wire tap_top0_pause_dr_o;
  wire tap_top0_update_dr_o;
  wire tap_top0_capture_dr_o;
  wire tap_top0_extest_select_o;
  wire tap_top0_sample_preload_select_o;
  wire tap_top0_mbist_select_o;
  wire tap_top0_debug_select_o;
  wire tap_top0_tdo_o;
  localparam n5759_o = 1'b0;
  localparam n5760_o = 1'b0;
  wire n5764_o;
  wire n5766_o;
  wire n5779_o;
  wire [1:0] n5780_o;
  wire n5783_o;
  wire n5786_o;
  wire [1:0] n5788_o;
  reg n5789_o;
  wire [1:0] n5791_o;
  wire [7:0] n5793_o;
  wire [63:0] n5794_o;
  wire [1:0] n5796_o;
  wire n5798_o;
  wire n5799_o;
  wire n5801_o;
  wire n5803_o;
  wire [72:0] n5805_o;
  wire [73:0] n5806_o;
  wire n5808_o;
  wire n5809_o;
  wire n5812_o;
  wire [1:0] n5814_o;
  wire [1:0] n5815_o;
  wire [1:0] n5816_o;
  wire [1:0] n5817_o;
  wire [71:0] n5818_o;
  wire [71:0] n5819_o;
  wire [71:0] n5820_o;
  wire n5821_o;
  wire n5822_o;
  wire n5823_o;
  wire [1:0] n5824_o;
  wire n5826_o;
  wire [63:0] n5827_o;
  wire [63:0] n5828_o;
  wire [63:0] n5829_o;
  wire [63:0] n5830_o;
  wire [63:0] n5831_o;
  wire [63:0] n5832_o;
  wire [63:0] n5833_o;
  wire [63:0] n5834_o;
  wire [7:0] n5835_o;
  wire [7:0] n5836_o;
  wire [7:0] n5837_o;
  wire [1:0] n5838_o;
  wire [1:0] n5839_o;
  wire [1:0] n5840_o;
  wire n5842_o;
  wire [71:0] n5843_o;
  wire [73:0] n5844_o;
  wire [73:0] n5845_o;
  wire [73:0] n5846_o;
  wire [73:0] n5848_o;
  wire [73:0] n5861_o;
  reg [73:0] n5862_q;
  wire [73:0] n5863_o;
  reg [73:0] n5864_q;
  wire n5865_o;
  reg n5866_q;
  reg n5867_q;
  reg n5868_q;
  reg n5869_q;
  reg n5870_q;
  assign dmi_addr = n5793_o;
  assign dmi_dout = n5794_o;
  assign dmi_req = jtag_req_1;
  assign dmi_wr = n5799_o;
  assign jtag_tdo = tap_top0_tdo_pad_o;
  /* dmi_dtm_jtag.vhdl:88:12  */
  assign capture = tap_top0_capture_dr_o; // (signal)
  /* dmi_dtm_jtag.vhdl:89:12  */
  assign update = tap_top0_update_dr_o; // (signal)
  /* dmi_dtm_jtag.vhdl:90:12  */
  assign sel = tap_top0_debug_select_o; // (signal)
  /* dmi_dtm_jtag.vhdl:91:12  */
  assign shift = tap_top0_shift_dr_o; // (signal)
  /* dmi_dtm_jtag.vhdl:92:12  */
  assign tdi = tap_top0_tdo_o; // (signal)
  /* dmi_dtm_jtag.vhdl:93:12  */
  assign tdo = n5801_o; // (signal)
  /* dmi_dtm_jtag.vhdl:98:12  */
  assign shiftr = n5862_q; // (signal)
  /* dmi_dtm_jtag.vhdl:101:12  */
  assign request = n5864_q; // (signal)
  /* dmi_dtm_jtag.vhdl:104:12  */
  assign jtag_req = n5866_q; // (signal)
  /* dmi_dtm_jtag.vhdl:107:12  */
  assign dmi_ack_0 = n5867_q; // (signal)
  /* dmi_dtm_jtag.vhdl:108:12  */
  assign dmi_ack_1 = n5868_q; // (signal)
  /* dmi_dtm_jtag.vhdl:113:12  */
  assign jtag_req_0 = n5869_q; // (signal)
  /* dmi_dtm_jtag.vhdl:114:12  */
  assign jtag_req_1 = n5870_q; // (signal)
  /* dmi_dtm_jtag.vhdl:117:12  */
  assign jtag_bsy = n5779_o; // (signal)
  /* dmi_dtm_jtag.vhdl:118:12  */
  assign op_valid = n5789_o; // (signal)
  /* dmi_dtm_jtag.vhdl:119:12  */
  assign rsp_op = n5791_o; // (signal)
  /* dmi_dtm_jtag.vhdl:166:5  */
  tap_top tap_top0 (
    .tms_pad_i(jtag_tms),
    .tck_pad_i(jtag_tck),
    .trst_pad_i(jtag_trst),
    .tdi_pad_i(jtag_tdi),
    .debug_tdi_i(tdo),
    .bs_chain_tdi_i(n5759_o),
    .mbist_tdi_i(n5760_o),
    .tdo_pad_o(tap_top0_tdo_pad_o),
    .tdo_padoe_o(),
    .shift_dr_o(tap_top0_shift_dr_o),
    .pause_dr_o(),
    .update_dr_o(tap_top0_update_dr_o),
    .capture_dr_o(tap_top0_capture_dr_o),
    .extest_select_o(),
    .sample_preload_select_o(),
    .mbist_select_o(),
    .debug_select_o(tap_top0_debug_select_o),
    .tdo_o(tap_top0_tdo_o));
  /* dmi_dtm_jtag.vhdl:197:13  */
  assign n5764_o = sys_reset ? 1'b0 : jtag_req;
  /* dmi_dtm_jtag.vhdl:197:13  */
  assign n5766_o = sys_reset ? 1'b0 : jtag_req_0;
  /* dmi_dtm_jtag.vhdl:225:26  */
  assign n5779_o = jtag_req | dmi_ack_1;
  /* dmi_dtm_jtag.vhdl:228:16  */
  assign n5780_o = shiftr[1:0];
  /* dmi_dtm_jtag.vhdl:229:13  */
  assign n5783_o = n5780_o == 2'b01;
  /* dmi_dtm_jtag.vhdl:230:13  */
  assign n5786_o = n5780_o == 2'b10;
  assign n5788_o = {n5786_o, n5783_o};
  /* dmi_dtm_jtag.vhdl:228:5  */
  always @*
    case (n5788_o)
      2'b10: n5789_o = 1'b1;
      2'b01: n5789_o = 1'b1;
      default: n5789_o = 1'b0;
    endcase
  /* dmi_dtm_jtag.vhdl:234:27  */
  assign n5791_o = jtag_bsy ? 2'b11 : 2'b00;
  /* dmi_dtm_jtag.vhdl:237:24  */
  assign n5793_o = request[73:66];
  /* dmi_dtm_jtag.vhdl:238:24  */
  assign n5794_o = request[65:2];
  /* dmi_dtm_jtag.vhdl:239:33  */
  assign n5796_o = request[1:0];
  /* dmi_dtm_jtag.vhdl:239:46  */
  assign n5798_o = n5796_o == 2'b10;
  /* dmi_dtm_jtag.vhdl:239:21  */
  assign n5799_o = n5798_o ? 1'b1 : 1'b0;
  /* dmi_dtm_jtag.vhdl:242:18  */
  assign n5801_o = shiftr[0];
  /* dmi_dtm_jtag.vhdl:250:28  */
  assign n5803_o = jtag_trst | sys_reset;
  /* dmi_dtm_jtag.vhdl:260:43  */
  assign n5805_o = shiftr[73:1];
  /* dmi_dtm_jtag.vhdl:260:35  */
  assign n5806_o = {tdi, n5805_o};
  /* dmi_dtm_jtag.vhdl:268:33  */
  assign n5808_o = update & op_valid;
  /* dmi_dtm_jtag.vhdl:269:33  */
  assign n5809_o = ~jtag_bsy;
  /* dmi_dtm_jtag.vhdl:268:17  */
  assign n5812_o = n5822_o ? 1'b1 : jtag_req;
  assign n5814_o = n5806_o[1:0];
  assign n5815_o = shiftr[1:0];
  /* dmi_dtm_jtag.vhdl:259:17  */
  assign n5816_o = shift ? n5814_o : n5815_o;
  /* dmi_dtm_jtag.vhdl:268:17  */
  assign n5817_o = n5808_o ? 2'b11 : n5816_o;
  assign n5818_o = n5806_o[73:2];
  assign n5819_o = shiftr[73:2];
  /* dmi_dtm_jtag.vhdl:259:17  */
  assign n5820_o = shift ? n5818_o : n5819_o;
  /* dmi_dtm_jtag.vhdl:268:17  */
  assign n5821_o = n5808_o & n5809_o;
  /* dmi_dtm_jtag.vhdl:268:17  */
  assign n5822_o = n5808_o & n5809_o;
  /* dmi_dtm_jtag.vhdl:287:35  */
  assign n5823_o = jtag_req & dmi_ack_1;
  /* dmi_dtm_jtag.vhdl:289:31  */
  assign n5824_o = request[1:0];
  /* dmi_dtm_jtag.vhdl:289:44  */
  assign n5826_o = n5824_o == 2'b01;
  assign n5827_o = shiftr[65:2];
  assign n5828_o = request[65:2];
  /* dmi_dtm_jtag.vhdl:268:17  */
  assign n5829_o = n5821_o ? n5827_o : n5828_o;
  /* dmi_dtm_jtag.vhdl:289:21  */
  assign n5830_o = n5826_o ? dmi_din : n5829_o;
  assign n5831_o = shiftr[65:2];
  assign n5832_o = request[65:2];
  /* dmi_dtm_jtag.vhdl:268:17  */
  assign n5833_o = n5821_o ? n5831_o : n5832_o;
  /* dmi_dtm_jtag.vhdl:287:17  */
  assign n5834_o = n5823_o ? n5830_o : n5833_o;
  assign n5835_o = shiftr[73:66];
  assign n5836_o = request[73:66];
  /* dmi_dtm_jtag.vhdl:268:17  */
  assign n5837_o = n5821_o ? n5835_o : n5836_o;
  assign n5838_o = shiftr[1:0];
  assign n5839_o = request[1:0];
  /* dmi_dtm_jtag.vhdl:268:17  */
  assign n5840_o = n5821_o ? n5838_o : n5839_o;
  /* dmi_dtm_jtag.vhdl:287:17  */
  assign n5842_o = n5823_o ? 1'b0 : n5812_o;
  /* dmi_dtm_jtag.vhdl:296:38  */
  assign n5843_o = request[73:2];
  /* dmi_dtm_jtag.vhdl:296:67  */
  assign n5844_o = {n5843_o, rsp_op};
  assign n5845_o = {n5820_o, n5817_o};
  /* dmi_dtm_jtag.vhdl:295:17  */
  assign n5846_o = capture ? n5844_o : n5845_o;
  assign n5848_o = {n5837_o, n5834_o, n5840_o};
  /* dmi_dtm_jtag.vhdl:254:9  */
  assign n5861_o = sel ? n5846_o : shiftr;
  /* dmi_dtm_jtag.vhdl:254:9  */
  always @(posedge jtag_tck or posedge n5803_o)
    if (n5803_o)
      n5862_q <= 74'b00000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n5862_q <= n5861_o;
  /* dmi_dtm_jtag.vhdl:254:9  */
  assign n5863_o = sel ? n5848_o : request;
  /* dmi_dtm_jtag.vhdl:254:9  */
  always @(posedge jtag_tck or posedge n5803_o)
    if (n5803_o)
      n5864_q <= 74'b00000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n5864_q <= n5863_o;
  /* dmi_dtm_jtag.vhdl:254:9  */
  assign n5865_o = sel ? n5842_o : jtag_req;
  /* dmi_dtm_jtag.vhdl:254:9  */
  always @(posedge jtag_tck or posedge n5803_o)
    if (n5803_o)
      n5866_q <= 1'b0;
    else
      n5866_q <= n5865_o;
  /* dmi_dtm_jtag.vhdl:215:9  */
  always @(posedge jtag_tck or posedge jtag_trst)
    if (jtag_trst)
      n5867_q <= 1'b0;
    else
      n5867_q <= dmi_ack;
  /* dmi_dtm_jtag.vhdl:215:9  */
  always @(posedge jtag_tck or posedge jtag_trst)
    if (jtag_trst)
      n5868_q <= 1'b0;
    else
      n5868_q <= dmi_ack_0;
  /* dmi_dtm_jtag.vhdl:196:9  */
  always @(posedge sys_clk)
    n5869_q <= n5764_o;
  /* dmi_dtm_jtag.vhdl:196:9  */
  always @(posedge sys_clk)
    n5870_q <= n5766_o;
endmodule

module wishbone_bram_wrapper_4096_a75adb9e07879fb6c63b494abe06e3f9a6bb2ed9
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  clk,
   input  rst,
   input  [28:0] wishbone_in_adr,
   input  [63:0] wishbone_in_dat,
   input  [7:0] wishbone_in_sel,
   input  wishbone_in_cyc,
   input  wishbone_in_stb,
   input  wishbone_in_we,
   output [63:0] wishbone_out_dat,
   output wishbone_out_ack,
   output wishbone_out_stall);
  wire [103:0] n5706_o;
  wire [63:0] n5708_o;
  wire n5709_o;
  wire n5710_o;
  wire [8:0] ram_addr;
  wire ram_we;
  wire ram_re;
  wire ack;
  wire ack_buf;
  wire [63:0] ram_0_dout;
  wire [63:0] n5711_o;
  wire [7:0] n5713_o;
  wire [8:0] n5714_o;
  wire n5715_o;
  wire n5716_o;
  wire n5717_o;
  wire n5718_o;
  wire n5719_o;
  wire n5720_o;
  wire n5721_o;
  wire n5722_o;
  wire n5723_o;
  wire n5724_o;
  wire n5725_o;
  wire n5729_o;
  wire n5730_o;
  wire n5731_o;
  wire n5732_o;
  wire n5733_o;
  wire n5734_o;
  wire n5735_o;
  wire n5737_o;
  wire n5739_o;
  wire n5741_o;
  reg n5745_q;
  reg n5746_q;
  wire [65:0] n5747_o;
  assign wishbone_out_dat = n5708_o;
  assign wishbone_out_ack = n5709_o;
  assign wishbone_out_stall = n5710_o;
  /* gpio.vhdl:25:9  */
  assign n5706_o = {wishbone_in_we, wishbone_in_stb, wishbone_in_cyc, wishbone_in_sel, wishbone_in_dat, wishbone_in_adr};
  /* gpio.vhdl:19:9  */
  assign n5708_o = n5747_o[63:0];
  assign n5709_o = n5747_o[64];
  /* gpio.vhdl:70:5  */
  assign n5710_o = n5747_o[65];
  /* wishbone_bram_wrapper.vhdl:30:12  */
  assign ram_addr = n5714_o; // (signal)
  /* wishbone_bram_wrapper.vhdl:31:12  */
  assign ram_we = n5719_o; // (signal)
  /* wishbone_bram_wrapper.vhdl:32:12  */
  assign ram_re = n5725_o; // (signal)
  /* wishbone_bram_wrapper.vhdl:35:12  */
  assign ack = n5745_q; // (signal)
  /* wishbone_bram_wrapper.vhdl:35:17  */
  assign ack_buf = n5746_q; // (signal)
  /* wishbone_bram_wrapper.vhdl:39:5  */
  main_bram_64_9_4096_a75adb9e07879fb6c63b494abe06e3f9a6bb2ed9 ram_0 (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(clk),
    .addr(ram_addr),
    .din(n5711_o),
    .sel(n5713_o),
    .re(ram_re),
    .we(ram_we),
    .dout(ram_0_dout));
  /* wishbone_bram_wrapper.vhdl:49:33  */
  assign n5711_o = n5706_o[92:29];
  /* wishbone_bram_wrapper.vhdl:51:32  */
  assign n5713_o = n5706_o[100:93];
  /* wishbone_bram_wrapper.vhdl:57:32  */
  assign n5714_o = n5706_o[8:0];
  /* wishbone_bram_wrapper.vhdl:58:27  */
  assign n5715_o = n5706_o[102];
  /* wishbone_bram_wrapper.vhdl:58:47  */
  assign n5716_o = n5706_o[101];
  /* wishbone_bram_wrapper.vhdl:58:31  */
  assign n5717_o = n5715_o & n5716_o;
  /* wishbone_bram_wrapper.vhdl:58:67  */
  assign n5718_o = n5706_o[103];
  /* wishbone_bram_wrapper.vhdl:58:51  */
  assign n5719_o = n5717_o & n5718_o;
  /* wishbone_bram_wrapper.vhdl:59:27  */
  assign n5720_o = n5706_o[102];
  /* wishbone_bram_wrapper.vhdl:59:47  */
  assign n5721_o = n5706_o[101];
  /* wishbone_bram_wrapper.vhdl:59:31  */
  assign n5722_o = n5720_o & n5721_o;
  /* wishbone_bram_wrapper.vhdl:59:71  */
  assign n5723_o = n5706_o[103];
  /* wishbone_bram_wrapper.vhdl:59:55  */
  assign n5724_o = ~n5723_o;
  /* wishbone_bram_wrapper.vhdl:59:51  */
  assign n5725_o = n5722_o & n5724_o;
  /* wishbone_bram_wrapper.vhdl:66:41  */
  assign n5729_o = n5706_o[101];
  /* wishbone_bram_wrapper.vhdl:66:45  */
  assign n5730_o = ~n5729_o;
  /* wishbone_bram_wrapper.vhdl:66:26  */
  assign n5731_o = rst | n5730_o;
  /* wishbone_bram_wrapper.vhdl:74:41  */
  assign n5732_o = ~ack;
  /* wishbone_bram_wrapper.vhdl:74:33  */
  assign n5733_o = ram_we & n5732_o;
  /* wishbone_bram_wrapper.vhdl:77:40  */
  assign n5734_o = n5706_o[102];
  /* wishbone_bram_wrapper.vhdl:74:17  */
  assign n5735_o = n5733_o ? ack : n5734_o;
  /* wishbone_bram_wrapper.vhdl:74:17  */
  assign n5737_o = n5733_o ? 1'b1 : ack;
  /* wishbone_bram_wrapper.vhdl:66:13  */
  assign n5739_o = n5731_o ? 1'b0 : n5735_o;
  /* wishbone_bram_wrapper.vhdl:66:13  */
  assign n5741_o = n5731_o ? 1'b0 : n5737_o;
  /* wishbone_bram_wrapper.vhdl:65:9  */
  always @(posedge clk)
    n5745_q <= n5739_o;
  /* wishbone_bram_wrapper.vhdl:65:9  */
  always @(posedge clk)
    n5746_q <= n5741_o;
  /* wishbone_bram_wrapper.vhdl:65:9  */
  assign n5747_o = {1'b0, ack_buf, ram_0_dout};
endmodule

module gpio_32
  (input  clk,
   input  rst,
   input  [29:0] wb_in_adr,
   input  [31:0] wb_in_dat,
   input  [3:0] wb_in_sel,
   input  wb_in_cyc,
   input  wb_in_stb,
   input  wb_in_we,
   input  [31:0] gpio_in,
   output [31:0] wb_out_dat,
   output wb_out_ack,
   output wb_out_stall,
   output [31:0] gpio_out,
   output [31:0] gpio_dir,
   output intr);
  wire [68:0] n5631_o;
  wire [31:0] n5633_o;
  wire n5634_o;
  wire n5635_o;
  reg [31:0] reg_data;
  reg [31:0] reg_dirn;
  wire [31:0] reg_in1;
  wire [31:0] reg_in2;
  wire [33:0] wb_rsp;
  wire [31:0] reg_out;
  localparam n5641_o = 1'b0;
  wire n5642_o;
  wire n5643_o;
  wire n5644_o;
  wire [4:0] n5645_o;
  wire n5647_o;
  wire n5649_o;
  wire n5651_o;
  wire [2:0] n5653_o;
  reg [31:0] n5654_o;
  wire n5659_o;
  wire n5660_o;
  wire n5661_o;
  wire n5662_o;
  wire n5663_o;
  wire [4:0] n5664_o;
  wire [31:0] n5665_o;
  wire n5667_o;
  wire [31:0] n5668_o;
  wire n5670_o;
  wire [31:0] n5671_o;
  wire [31:0] n5672_o;
  wire n5674_o;
  wire [31:0] n5675_o;
  wire [31:0] n5676_o;
  wire [31:0] n5677_o;
  wire n5679_o;
  wire [3:0] n5680_o;
  reg [31:0] n5681_o;
  reg [31:0] n5682_o;
  wire [31:0] n5683_o;
  wire [31:0] n5684_o;
  wire n5685_o;
  wire n5686_o;
  wire n5687_o;
  wire [31:0] n5688_o;
  wire [31:0] n5690_o;
  wire [31:0] n5692_o;
  wire [33:0] n5693_o;
  reg [31:0] n5700_q;
  reg [31:0] n5701_q;
  reg [31:0] n5702_q;
  reg [31:0] n5703_q;
  wire [33:0] n5704_o;
  reg [33:0] n5705_q;
  assign wb_out_dat = n5633_o;
  assign wb_out_ack = n5634_o;
  assign wb_out_stall = n5635_o;
  assign gpio_out = reg_data;
  assign gpio_dir = reg_dirn;
  assign intr = n5641_o;
  /* xics.vhdl:295:9  */
  assign n5631_o = {wb_in_we, wb_in_stb, wb_in_cyc, wb_in_sel, wb_in_dat, wb_in_adr};
  assign n5633_o = n5705_q[31:0];
  assign n5634_o = n5705_q[32];
  assign n5635_o = n5705_q[33];
  /* gpio.vhdl:43:12  */
  always @*
    reg_data = n5700_q; // (isignal)
  initial
    reg_data = 32'b00000000000000000000000000000000;
  /* gpio.vhdl:44:12  */
  always @*
    reg_dirn = n5701_q; // (isignal)
  initial
    reg_dirn = 32'b00000000000000000000000000000000;
  /* gpio.vhdl:45:12  */
  assign reg_in1 = n5702_q; // (signal)
  /* gpio.vhdl:46:12  */
  assign reg_in2 = n5703_q; // (signal)
  /* gpio.vhdl:48:12  */
  assign wb_rsp = n5704_o; // (signal)
  /* gpio.vhdl:49:12  */
  assign reg_out = n5654_o; // (signal)
  /* gpio.vhdl:60:25  */
  assign n5642_o = n5631_o[66];
  /* gpio.vhdl:60:39  */
  assign n5643_o = n5631_o[67];
  /* gpio.vhdl:60:29  */
  assign n5644_o = n5642_o & n5643_o;
  /* gpio.vhdl:61:19  */
  assign n5645_o = n5631_o[4:0];
  /* gpio.vhdl:62:18  */
  assign n5647_o = n5645_o == 5'b00000;
  /* gpio.vhdl:63:18  */
  assign n5649_o = n5645_o == 5'b00001;
  /* gpio.vhdl:64:18  */
  assign n5651_o = n5645_o == 5'b00010;
  assign n5653_o = {n5651_o, n5649_o, n5647_o};
  /* gpio.vhdl:61:5  */
  always @*
    case (n5653_o)
      3'b100: n5654_o = reg_dirn;
      3'b010: n5654_o = reg_in2;
      3'b001: n5654_o = reg_data;
      default: n5654_o = 32'b00000000000000000000000000000000;
    endcase
  /* gpio.vhdl:81:26  */
  assign n5659_o = n5631_o[66];
  /* gpio.vhdl:81:46  */
  assign n5660_o = n5631_o[67];
  /* gpio.vhdl:81:36  */
  assign n5661_o = n5659_o & n5660_o;
  /* gpio.vhdl:81:66  */
  assign n5662_o = n5631_o[68];
  /* gpio.vhdl:81:56  */
  assign n5663_o = n5661_o & n5662_o;
  /* gpio.vhdl:82:35  */
  assign n5664_o = n5631_o[4:0];
  /* gpio.vhdl:84:50  */
  assign n5665_o = n5631_o[61:30];
  /* gpio.vhdl:83:25  */
  assign n5667_o = n5664_o == 5'b00000;
  /* gpio.vhdl:86:50  */
  assign n5668_o = n5631_o[61:30];
  /* gpio.vhdl:85:25  */
  assign n5670_o = n5664_o == 5'b00010;
  /* gpio.vhdl:88:62  */
  assign n5671_o = n5631_o[61:30];
  /* gpio.vhdl:88:50  */
  assign n5672_o = reg_data | n5671_o;
  /* gpio.vhdl:87:25  */
  assign n5674_o = n5664_o == 5'b00100;
  /* gpio.vhdl:90:67  */
  assign n5675_o = n5631_o[61:30];
  /* gpio.vhdl:90:54  */
  assign n5676_o = ~n5675_o;
  /* gpio.vhdl:90:50  */
  assign n5677_o = reg_data & n5676_o;
  /* gpio.vhdl:89:25  */
  assign n5679_o = n5664_o == 5'b00101;
  assign n5680_o = {n5679_o, n5674_o, n5670_o, n5667_o};
  /* gpio.vhdl:82:21  */
  always @*
    case (n5680_o)
      4'b1000: n5681_o = n5677_o;
      4'b0100: n5681_o = n5672_o;
      4'b0010: n5681_o = reg_data;
      4'b0001: n5681_o = n5665_o;
      default: n5681_o = reg_data;
    endcase
  /* gpio.vhdl:82:21  */
  always @*
    case (n5680_o)
      4'b1000: n5682_o = reg_dirn;
      4'b0100: n5682_o = reg_dirn;
      4'b0010: n5682_o = n5668_o;
      4'b0001: n5682_o = reg_dirn;
      default: n5682_o = reg_dirn;
    endcase
  /* gpio.vhdl:81:17  */
  assign n5683_o = n5663_o ? n5681_o : reg_data;
  /* gpio.vhdl:81:17  */
  assign n5684_o = n5663_o ? n5682_o : reg_dirn;
  assign n5685_o = wb_rsp[32];
  /* gpio.vhdl:76:13  */
  assign n5686_o = rst ? 1'b0 : n5685_o;
  assign n5687_o = wb_rsp[33];
  assign n5688_o = wb_rsp[31:0];
  /* gpio.vhdl:76:13  */
  assign n5690_o = rst ? 32'b00000000000000000000000000000000 : n5683_o;
  /* gpio.vhdl:76:13  */
  assign n5692_o = rst ? 32'b00000000000000000000000000000000 : n5684_o;
  assign n5693_o = {n5687_o, n5686_o, n5688_o};
  /* gpio.vhdl:72:9  */
  always @(posedge clk)
    n5700_q <= n5690_o;
  initial
    n5700_q = 32'b00000000000000000000000000000000;
  /* gpio.vhdl:72:9  */
  always @(posedge clk)
    n5701_q <= n5692_o;
  initial
    n5701_q = 32'b00000000000000000000000000000000;
  /* gpio.vhdl:72:9  */
  always @(posedge clk)
    n5702_q <= gpio_in;
  /* gpio.vhdl:72:9  */
  always @(posedge clk)
    n5703_q <= reg_in1;
  /* gpio.vhdl:72:9  */
  assign n5704_o = {1'b0, n5644_o, reg_out};
  /* gpio.vhdl:72:9  */
  always @(posedge clk)
    n5705_q <= n5693_o;
endmodule

module xics_ics_16_3
  (input  clk,
   input  rst,
   input  [29:0] wb_in_adr,
   input  [31:0] wb_in_dat,
   input  [3:0] wb_in_sel,
   input  wb_in_cyc,
   input  wb_in_stb,
   input  wb_in_we,
   input  [15:0] int_level_in,
   output [31:0] wb_out_dat,
   output wb_out_ack,
   output wb_out_stall,
   output [3:0] icp_out_src,
   output [7:0] icp_out_pri);
  wire [68:0] n3081_o;
  wire [31:0] n3083_o;
  wire n3084_o;
  wire n3085_o;
  wire [3:0] n3087_o;
  wire [7:0] n3088_o;
  wire [47:0] xives;
  wire wb_valid;
  wire [3:0] reg_idx;
  wire [11:0] icp_out_next;
  wire [15:0] int_level_l;
  wire reg_is_xive;
  wire reg_is_config;
  wire reg_is_debug;
  wire n3089_o;
  wire [9:0] n3091_o;
  wire n3093_o;
  wire n3094_o;
  wire [9:0] n3097_o;
  wire n3099_o;
  wire n3100_o;
  wire [3:0] n3102_o;
  wire n3109_o;
  wire n3110_o;
  wire n3111_o;
  wire [1:0] n3118_o;
  wire [2:0] n3121_o;
  wire [3:0] n3123_o;
  wire [23:0] n3125_o;
  wire [3:0] n3128_o;
  wire [2:0] n3131_o;
  wire n3138_o;
  localparam [7:0] n3139_o = 8'b00000000;
  wire [4:0] n3140_o;
  wire [7:0] n3141_o;
  wire [7:0] n3143_o;
  wire [31:0] n3145_o;
  wire [3:0] n3147_o;
  wire [23:0] n3149_o;
  wire [7:0] n3150_o;
  wire [31:0] n3151_o;
  wire [31:0] n3153_o;
  wire [31:0] n3155_o;
  wire [31:0] n3156_o;
  wire [7:0] n3164_o;
  wire [7:0] n3167_o;
  wire [7:0] n3169_o;
  wire [7:0] n3171_o;
  wire [31:0] n3172_o;
  wire [32:0] n3173_o;
  wire [31:0] n3181_o;
  wire [7:0] n3187_o;
  wire [7:0] n3190_o;
  wire [7:0] n3192_o;
  wire [7:0] n3194_o;
  wire [31:0] n3195_o;
  wire n3213_o;
  wire n3214_o;
  wire [3:0] n3216_o;
  wire [7:0] n3219_o;
  localparam [7:0] n3226_o = 8'b00000000;
  wire [4:0] n3227_o;
  wire [7:0] n3228_o;
  wire n3229_o;
  wire [2:0] n3231_o;
  wire [2:0] n3232_o;
  wire [47:0] n3234_o;
  wire n3235_o;
  wire [47:0] n3236_o;
  wire [47:0] n3237_o;
  wire n3249_o;
  wire [2:0] n3251_o;
  wire [2:0] n3252_o;
  localparam [7:0] n3260_o = 8'b00000000;
  wire [7:0] n3265_o;
  localparam [7:0] n3266_o = 8'b00000000;
  wire [7:0] n3267_o;
  wire n3269_o;
  wire [2:0] n3271_o;
  wire [2:0] n3272_o;
  localparam [7:0] n3280_o = 8'b00000000;
  wire [7:0] n3284_o;
  wire [7:0] n3285_o;
  wire n3286_o;
  wire [2:0] n3288_o;
  wire [2:0] n3289_o;
  localparam [7:0] n3297_o = 8'b00000000;
  wire [7:0] n3301_o;
  wire [7:0] n3302_o;
  wire n3303_o;
  wire [2:0] n3305_o;
  wire [2:0] n3306_o;
  localparam [7:0] n3314_o = 8'b00000000;
  wire [7:0] n3318_o;
  wire [7:0] n3319_o;
  wire n3320_o;
  wire [2:0] n3322_o;
  wire [2:0] n3323_o;
  localparam [7:0] n3331_o = 8'b00000000;
  wire [7:0] n3335_o;
  wire [7:0] n3336_o;
  wire n3337_o;
  wire [2:0] n3339_o;
  wire [2:0] n3340_o;
  localparam [7:0] n3348_o = 8'b00000000;
  wire [7:0] n3352_o;
  wire [7:0] n3353_o;
  wire n3354_o;
  wire [2:0] n3356_o;
  wire [2:0] n3357_o;
  localparam [7:0] n3365_o = 8'b00000000;
  wire [7:0] n3369_o;
  wire [7:0] n3370_o;
  wire n3371_o;
  wire [2:0] n3373_o;
  wire [2:0] n3374_o;
  localparam [7:0] n3382_o = 8'b00000000;
  wire [7:0] n3386_o;
  wire [7:0] n3387_o;
  wire n3388_o;
  wire [2:0] n3390_o;
  wire [2:0] n3391_o;
  localparam [7:0] n3399_o = 8'b00000000;
  wire [7:0] n3403_o;
  wire [7:0] n3404_o;
  wire n3405_o;
  wire [2:0] n3407_o;
  wire [2:0] n3408_o;
  localparam [7:0] n3416_o = 8'b00000000;
  wire [7:0] n3420_o;
  wire [7:0] n3421_o;
  wire n3422_o;
  wire [2:0] n3424_o;
  wire [2:0] n3425_o;
  localparam [7:0] n3433_o = 8'b00000000;
  wire [7:0] n3437_o;
  wire [7:0] n3438_o;
  wire n3439_o;
  wire [2:0] n3441_o;
  wire [2:0] n3442_o;
  localparam [7:0] n3450_o = 8'b00000000;
  wire [7:0] n3454_o;
  wire [7:0] n3455_o;
  wire n3456_o;
  wire [2:0] n3458_o;
  wire [2:0] n3459_o;
  localparam [7:0] n3467_o = 8'b00000000;
  wire [7:0] n3471_o;
  wire [7:0] n3472_o;
  wire n3473_o;
  wire [2:0] n3475_o;
  wire [2:0] n3476_o;
  localparam [7:0] n3484_o = 8'b00000000;
  wire [7:0] n3488_o;
  wire [7:0] n3489_o;
  wire n3490_o;
  wire [2:0] n3492_o;
  wire [2:0] n3493_o;
  localparam [7:0] n3501_o = 8'b00000000;
  wire [7:0] n3505_o;
  wire [7:0] n3506_o;
  wire n3507_o;
  wire [2:0] n3509_o;
  wire [2:0] n3510_o;
  localparam [7:0] n3518_o = 8'b00000000;
  wire [7:0] n3522_o;
  wire [6:0] n3533_o;
  wire [6:0] n3534_o;
  wire [6:0] n3535_o;
  wire [6:0] n3536_o;
  wire [6:0] n3537_o;
  wire [6:0] n3538_o;
  wire [6:0] n3539_o;
  wire [6:0] n3540_o;
  wire [6:0] n3541_o;
  wire [6:0] n3542_o;
  wire [6:0] n3543_o;
  wire [6:0] n3544_o;
  wire [6:0] n3545_o;
  wire [6:0] n3546_o;
  wire [6:0] n3547_o;
  wire [6:0] n3548_o;
  wire [6:0] n3549_o;
  wire [6:0] n3550_o;
  wire [6:0] n3551_o;
  wire [6:0] n3552_o;
  wire [6:0] n3553_o;
  wire [6:0] n3554_o;
  wire [6:0] n3555_o;
  wire [6:0] n3556_o;
  wire [6:0] n3557_o;
  wire [6:0] n3558_o;
  wire [6:0] n3559_o;
  wire [6:0] n3560_o;
  wire [6:0] n3561_o;
  wire [6:0] n3562_o;
  wire [6:0] n3563_o;
  wire [6:0] n3564_o;
  wire [6:0] n3565_o;
  wire [7:0] n3577_o;
  wire [7:0] n3578_o;
  wire [7:0] n3580_o;
  wire [7:0] n3581_o;
  wire [7:0] n3583_o;
  wire [7:0] n3584_o;
  wire [63:0] n3587_o;
  wire n3596_o;
  wire n3597_o;
  wire n3598_o;
  wire n3599_o;
  wire n3601_o;
  wire n3603_o;
  wire n3604_o;
  wire n3605_o;
  wire n3606_o;
  wire n3607_o;
  wire n3608_o;
  wire n3609_o;
  wire n3610_o;
  wire n3611_o;
  wire n3612_o;
  wire n3613_o;
  wire n3614_o;
  wire n3615_o;
  wire n3616_o;
  wire n3617_o;
  wire n3618_o;
  wire n3619_o;
  wire n3620_o;
  wire n3621_o;
  wire n3622_o;
  wire n3623_o;
  wire n3624_o;
  wire n3625_o;
  wire n3626_o;
  wire n3627_o;
  wire n3628_o;
  wire n3629_o;
  wire n3630_o;
  wire n3631_o;
  wire n3632_o;
  wire n3633_o;
  wire n3634_o;
  wire n3635_o;
  wire n3636_o;
  wire n3637_o;
  wire n3638_o;
  wire n3639_o;
  wire n3640_o;
  wire n3641_o;
  wire n3642_o;
  wire n3643_o;
  wire n3644_o;
  wire n3645_o;
  wire n3646_o;
  wire n3647_o;
  wire n3648_o;
  wire n3649_o;
  wire n3650_o;
  wire n3651_o;
  wire n3652_o;
  wire n3653_o;
  wire n3654_o;
  wire n3655_o;
  wire n3656_o;
  wire n3657_o;
  wire n3658_o;
  wire n3659_o;
  wire n3660_o;
  wire n3661_o;
  wire n3662_o;
  wire n3663_o;
  wire n3664_o;
  wire n3665_o;
  wire n3666_o;
  wire n3667_o;
  wire n3668_o;
  wire n3669_o;
  wire n3670_o;
  wire n3671_o;
  wire n3672_o;
  wire n3673_o;
  wire n3674_o;
  wire n3675_o;
  wire n3676_o;
  wire n3677_o;
  wire n3678_o;
  wire n3679_o;
  wire n3680_o;
  wire n3681_o;
  wire n3682_o;
  wire n3683_o;
  wire n3684_o;
  wire n3685_o;
  wire n3686_o;
  wire n3687_o;
  wire n3688_o;
  wire n3689_o;
  wire n3690_o;
  wire n3691_o;
  wire n3692_o;
  wire n3693_o;
  wire n3694_o;
  wire n3695_o;
  wire n3696_o;
  wire n3697_o;
  wire n3698_o;
  wire n3699_o;
  wire n3700_o;
  wire n3701_o;
  wire n3702_o;
  wire n3703_o;
  wire n3704_o;
  wire n3705_o;
  wire n3706_o;
  wire n3707_o;
  wire n3708_o;
  wire n3709_o;
  wire n3710_o;
  wire n3711_o;
  wire n3712_o;
  wire n3713_o;
  wire n3714_o;
  wire n3715_o;
  wire n3716_o;
  wire n3717_o;
  wire n3718_o;
  wire n3719_o;
  wire n3720_o;
  wire n3721_o;
  wire n3722_o;
  wire n3723_o;
  wire n3724_o;
  wire n3725_o;
  wire n3726_o;
  wire n3727_o;
  wire n3728_o;
  wire n3729_o;
  wire n3730_o;
  wire n3731_o;
  wire n3732_o;
  wire n3733_o;
  wire n3734_o;
  wire n3735_o;
  wire n3736_o;
  wire n3737_o;
  wire n3738_o;
  wire n3739_o;
  wire n3740_o;
  wire n3741_o;
  wire n3742_o;
  wire n3743_o;
  wire n3744_o;
  wire n3745_o;
  wire n3746_o;
  wire n3747_o;
  wire n3748_o;
  wire n3749_o;
  wire n3750_o;
  wire n3751_o;
  wire n3752_o;
  wire n3753_o;
  wire n3754_o;
  wire n3755_o;
  wire n3756_o;
  wire n3757_o;
  wire n3760_o;
  wire n3761_o;
  wire n3762_o;
  wire n3763_o;
  wire n3765_o;
  wire n3767_o;
  wire n3768_o;
  wire n3769_o;
  wire n3770_o;
  wire n3771_o;
  wire n3772_o;
  wire n3773_o;
  wire n3774_o;
  wire n3775_o;
  wire n3776_o;
  wire n3777_o;
  wire n3778_o;
  wire n3779_o;
  wire n3780_o;
  wire n3781_o;
  wire n3782_o;
  wire n3783_o;
  wire n3784_o;
  wire n3785_o;
  wire n3786_o;
  wire n3787_o;
  wire n3788_o;
  wire n3789_o;
  wire n3790_o;
  wire n3791_o;
  wire n3792_o;
  wire n3793_o;
  wire n3794_o;
  wire n3795_o;
  wire n3796_o;
  wire n3797_o;
  wire n3798_o;
  wire n3799_o;
  wire n3800_o;
  wire n3801_o;
  wire n3802_o;
  wire n3803_o;
  wire n3804_o;
  wire n3805_o;
  wire n3806_o;
  wire n3807_o;
  wire n3808_o;
  wire n3809_o;
  wire n3810_o;
  wire n3811_o;
  wire n3812_o;
  wire n3813_o;
  wire n3814_o;
  wire n3815_o;
  wire n3816_o;
  wire n3817_o;
  wire n3818_o;
  wire n3819_o;
  wire n3820_o;
  wire n3821_o;
  wire n3822_o;
  wire n3823_o;
  wire n3824_o;
  wire n3825_o;
  wire n3826_o;
  wire n3827_o;
  wire n3828_o;
  wire n3829_o;
  wire n3830_o;
  wire n3831_o;
  wire n3832_o;
  wire n3833_o;
  wire n3834_o;
  wire n3835_o;
  wire n3836_o;
  wire n3837_o;
  wire n3838_o;
  wire n3839_o;
  wire n3840_o;
  wire n3841_o;
  wire n3843_o;
  wire n3844_o;
  wire n3845_o;
  wire n3846_o;
  wire n3848_o;
  wire n3850_o;
  wire n3851_o;
  wire n3852_o;
  wire n3853_o;
  wire n3854_o;
  wire n3855_o;
  wire n3856_o;
  wire n3857_o;
  wire n3858_o;
  wire n3859_o;
  wire n3860_o;
  wire n3861_o;
  wire n3862_o;
  wire n3863_o;
  wire n3864_o;
  wire n3865_o;
  wire n3866_o;
  wire n3867_o;
  wire n3868_o;
  wire n3869_o;
  wire n3870_o;
  wire n3871_o;
  wire n3872_o;
  wire n3873_o;
  wire n3874_o;
  wire n3875_o;
  wire n3876_o;
  wire n3877_o;
  wire n3878_o;
  wire n3879_o;
  wire n3880_o;
  wire n3881_o;
  wire n3882_o;
  wire n3883_o;
  wire n3884_o;
  wire n3886_o;
  wire n3887_o;
  wire n3888_o;
  wire n3889_o;
  wire n3891_o;
  wire n3893_o;
  wire n3894_o;
  wire n3895_o;
  wire n3896_o;
  wire n3897_o;
  wire n3898_o;
  wire n3899_o;
  wire n3900_o;
  wire n3901_o;
  wire n3902_o;
  wire n3903_o;
  wire n3904_o;
  wire n3905_o;
  wire n3906_o;
  wire n3907_o;
  wire n3909_o;
  wire n3910_o;
  wire n3911_o;
  wire n3912_o;
  wire n3914_o;
  wire n3916_o;
  wire n3917_o;
  wire n3918_o;
  wire n3919_o;
  wire n3920_o;
  wire n3922_o;
  wire n3923_o;
  wire n3924_o;
  wire n3925_o;
  wire n3927_o;
  wire [5:0] n3929_o;
  wire [63:0] n3932_o;
  wire n3941_o;
  wire n3942_o;
  wire n3944_o;
  wire n3946_o;
  wire n3947_o;
  wire n3948_o;
  wire n3949_o;
  wire n3950_o;
  wire n3951_o;
  wire n3952_o;
  wire n3953_o;
  wire n3954_o;
  wire n3955_o;
  wire n3956_o;
  wire n3957_o;
  wire n3958_o;
  wire n3959_o;
  wire n3960_o;
  wire n3961_o;
  wire n3962_o;
  wire n3963_o;
  wire n3964_o;
  wire n3965_o;
  wire n3966_o;
  wire n3967_o;
  wire n3968_o;
  wire n3969_o;
  wire n3970_o;
  wire n3971_o;
  wire n3972_o;
  wire n3973_o;
  wire n3974_o;
  wire n3975_o;
  wire n3976_o;
  wire n3977_o;
  wire n3978_o;
  wire n3979_o;
  wire n3980_o;
  wire n3981_o;
  wire n3982_o;
  wire n3983_o;
  wire n3984_o;
  wire n3985_o;
  wire n3986_o;
  wire n3987_o;
  wire n3988_o;
  wire n3989_o;
  wire n3990_o;
  wire n3991_o;
  wire n3992_o;
  wire n3993_o;
  wire n3994_o;
  wire n3995_o;
  wire n3996_o;
  wire n3997_o;
  wire n3998_o;
  wire n3999_o;
  wire n4000_o;
  wire n4001_o;
  wire n4002_o;
  wire n4003_o;
  wire n4004_o;
  wire n4005_o;
  wire n4006_o;
  wire n4007_o;
  wire n4008_o;
  wire n4009_o;
  wire n4010_o;
  wire n4011_o;
  wire n4012_o;
  wire n4013_o;
  wire n4014_o;
  wire n4015_o;
  wire n4016_o;
  wire n4017_o;
  wire n4018_o;
  wire n4019_o;
  wire n4020_o;
  wire n4021_o;
  wire n4022_o;
  wire n4023_o;
  wire n4024_o;
  wire n4025_o;
  wire n4026_o;
  wire n4027_o;
  wire n4028_o;
  wire n4029_o;
  wire n4030_o;
  wire n4031_o;
  wire n4032_o;
  wire n4033_o;
  wire n4034_o;
  wire n4035_o;
  wire n4036_o;
  wire n4037_o;
  wire n4038_o;
  wire [1:0] n4041_o;
  wire n4042_o;
  wire n4044_o;
  wire [1:0] n4046_o;
  wire n4047_o;
  wire n4048_o;
  wire [1:0] n4049_o;
  wire n4050_o;
  wire n4051_o;
  wire [1:0] n4052_o;
  wire n4053_o;
  wire n4054_o;
  wire [1:0] n4055_o;
  wire n4056_o;
  wire n4057_o;
  wire [1:0] n4058_o;
  wire n4059_o;
  wire n4060_o;
  wire [1:0] n4061_o;
  wire n4062_o;
  wire n4063_o;
  wire [1:0] n4064_o;
  wire n4065_o;
  wire n4066_o;
  wire [1:0] n4067_o;
  wire n4068_o;
  wire n4069_o;
  wire [1:0] n4070_o;
  wire n4071_o;
  wire n4072_o;
  wire [1:0] n4073_o;
  wire n4074_o;
  wire n4075_o;
  wire [1:0] n4076_o;
  wire n4077_o;
  wire n4078_o;
  wire [1:0] n4079_o;
  wire n4080_o;
  wire n4081_o;
  wire [1:0] n4082_o;
  wire n4083_o;
  wire n4084_o;
  wire [1:0] n4085_o;
  wire n4086_o;
  wire n4087_o;
  wire [1:0] n4088_o;
  wire n4089_o;
  wire n4090_o;
  wire [3:0] n4092_o;
  wire n4093_o;
  wire n4095_o;
  wire [3:0] n4097_o;
  wire n4098_o;
  wire n4099_o;
  wire [3:0] n4100_o;
  wire n4101_o;
  wire n4102_o;
  wire [3:0] n4103_o;
  wire n4104_o;
  wire n4105_o;
  wire [3:0] n4106_o;
  wire n4107_o;
  wire n4108_o;
  wire [3:0] n4109_o;
  wire n4110_o;
  wire n4111_o;
  wire [3:0] n4112_o;
  wire n4113_o;
  wire n4114_o;
  wire [3:0] n4115_o;
  wire n4116_o;
  wire n4117_o;
  wire [7:0] n4119_o;
  wire n4120_o;
  wire n4122_o;
  wire [7:0] n4124_o;
  wire n4125_o;
  wire n4126_o;
  wire [7:0] n4127_o;
  wire n4128_o;
  wire n4129_o;
  wire [7:0] n4130_o;
  wire n4131_o;
  wire n4132_o;
  wire [15:0] n4134_o;
  wire n4135_o;
  wire n4137_o;
  wire [15:0] n4139_o;
  wire n4140_o;
  wire n4141_o;
  wire [31:0] n4143_o;
  wire n4144_o;
  wire n4146_o;
  wire [5:0] n4148_o;
  wire [3:0] n4150_o;
  wire [1:0] n4151_o;
  wire [5:0] n4152_o;
  wire [2:0] n4155_o;
  wire n4156_o;
  wire [2:0] n4157_o;
  wire [2:0] n4158_o;
  wire n4159_o;
  wire n4160_o;
  wire n4163_o;
  localparam [15:0] n4164_o = 16'b0000000000000000;
  wire n4166_o;
  wire [2:0] n4167_o;
  wire [2:0] n4168_o;
  wire n4169_o;
  wire n4170_o;
  wire n4172_o;
  wire n4173_o;
  wire n4175_o;
  wire [2:0] n4176_o;
  wire [2:0] n4177_o;
  wire n4178_o;
  wire n4179_o;
  wire n4181_o;
  wire n4182_o;
  wire n4184_o;
  wire [2:0] n4185_o;
  wire [2:0] n4186_o;
  wire n4187_o;
  wire n4188_o;
  wire n4190_o;
  wire n4191_o;
  wire n4193_o;
  wire [2:0] n4194_o;
  wire [2:0] n4195_o;
  wire n4196_o;
  wire n4197_o;
  wire n4199_o;
  wire n4200_o;
  wire n4202_o;
  wire [2:0] n4203_o;
  wire [2:0] n4204_o;
  wire n4205_o;
  wire n4206_o;
  wire n4208_o;
  wire n4209_o;
  wire n4211_o;
  wire [2:0] n4212_o;
  wire [2:0] n4213_o;
  wire n4214_o;
  wire n4215_o;
  wire n4217_o;
  wire n4218_o;
  wire n4220_o;
  wire [2:0] n4221_o;
  wire [2:0] n4222_o;
  wire n4223_o;
  wire n4224_o;
  wire n4226_o;
  wire n4227_o;
  wire n4229_o;
  wire [2:0] n4230_o;
  wire [2:0] n4231_o;
  wire n4232_o;
  wire n4233_o;
  wire n4235_o;
  wire n4236_o;
  wire n4238_o;
  wire [2:0] n4239_o;
  wire [2:0] n4240_o;
  wire n4241_o;
  wire n4242_o;
  wire n4244_o;
  wire n4245_o;
  wire n4247_o;
  wire [2:0] n4248_o;
  wire [2:0] n4249_o;
  wire n4250_o;
  wire n4251_o;
  wire n4253_o;
  wire n4254_o;
  wire n4256_o;
  wire [2:0] n4257_o;
  wire [2:0] n4258_o;
  wire n4259_o;
  wire n4260_o;
  wire n4262_o;
  wire n4263_o;
  wire n4265_o;
  wire [2:0] n4266_o;
  wire [2:0] n4267_o;
  wire n4268_o;
  wire n4269_o;
  wire n4271_o;
  wire n4272_o;
  wire n4274_o;
  wire [2:0] n4275_o;
  wire [2:0] n4276_o;
  wire n4277_o;
  wire n4278_o;
  wire n4280_o;
  wire n4281_o;
  wire n4283_o;
  wire [2:0] n4284_o;
  wire [2:0] n4285_o;
  wire n4286_o;
  wire n4287_o;
  wire n4289_o;
  wire n4290_o;
  wire n4291_o;
  wire n4292_o;
  wire [2:0] n4293_o;
  wire [2:0] n4294_o;
  wire n4295_o;
  wire n4296_o;
  wire n4298_o;
  wire [15:0] n4306_o;
  wire [14:0] n4309_o;
  wire [15:0] n4321_o;
  wire [15:0] n4322_o;
  wire [15:0] n4324_o;
  wire [15:0] n4325_o;
  wire [15:0] n4327_o;
  wire [15:0] n4328_o;
  wire [63:0] n4331_o;
  wire n4340_o;
  wire n4341_o;
  wire n4342_o;
  wire n4343_o;
  wire n4345_o;
  wire n4347_o;
  wire n4348_o;
  wire n4349_o;
  wire n4350_o;
  wire n4351_o;
  wire n4352_o;
  wire n4353_o;
  wire n4354_o;
  wire n4355_o;
  wire n4356_o;
  wire n4357_o;
  wire n4358_o;
  wire n4359_o;
  wire n4360_o;
  wire n4361_o;
  wire n4362_o;
  wire n4363_o;
  wire n4364_o;
  wire n4365_o;
  wire n4366_o;
  wire n4367_o;
  wire n4368_o;
  wire n4369_o;
  wire n4370_o;
  wire n4371_o;
  wire n4372_o;
  wire n4373_o;
  wire n4374_o;
  wire n4375_o;
  wire n4376_o;
  wire n4377_o;
  wire n4378_o;
  wire n4379_o;
  wire n4380_o;
  wire n4381_o;
  wire n4382_o;
  wire n4383_o;
  wire n4384_o;
  wire n4385_o;
  wire n4386_o;
  wire n4387_o;
  wire n4388_o;
  wire n4389_o;
  wire n4390_o;
  wire n4391_o;
  wire n4392_o;
  wire n4393_o;
  wire n4394_o;
  wire n4395_o;
  wire n4396_o;
  wire n4397_o;
  wire n4398_o;
  wire n4399_o;
  wire n4400_o;
  wire n4401_o;
  wire n4402_o;
  wire n4403_o;
  wire n4404_o;
  wire n4405_o;
  wire n4406_o;
  wire n4407_o;
  wire n4408_o;
  wire n4409_o;
  wire n4410_o;
  wire n4411_o;
  wire n4412_o;
  wire n4413_o;
  wire n4414_o;
  wire n4415_o;
  wire n4416_o;
  wire n4417_o;
  wire n4418_o;
  wire n4419_o;
  wire n4420_o;
  wire n4421_o;
  wire n4422_o;
  wire n4423_o;
  wire n4424_o;
  wire n4425_o;
  wire n4426_o;
  wire n4427_o;
  wire n4428_o;
  wire n4429_o;
  wire n4430_o;
  wire n4431_o;
  wire n4432_o;
  wire n4433_o;
  wire n4434_o;
  wire n4435_o;
  wire n4436_o;
  wire n4437_o;
  wire n4438_o;
  wire n4439_o;
  wire n4440_o;
  wire n4441_o;
  wire n4442_o;
  wire n4443_o;
  wire n4444_o;
  wire n4445_o;
  wire n4446_o;
  wire n4447_o;
  wire n4448_o;
  wire n4449_o;
  wire n4450_o;
  wire n4451_o;
  wire n4452_o;
  wire n4453_o;
  wire n4454_o;
  wire n4455_o;
  wire n4456_o;
  wire n4457_o;
  wire n4458_o;
  wire n4459_o;
  wire n4460_o;
  wire n4461_o;
  wire n4462_o;
  wire n4463_o;
  wire n4464_o;
  wire n4465_o;
  wire n4466_o;
  wire n4467_o;
  wire n4468_o;
  wire n4469_o;
  wire n4470_o;
  wire n4471_o;
  wire n4472_o;
  wire n4473_o;
  wire n4474_o;
  wire n4475_o;
  wire n4476_o;
  wire n4477_o;
  wire n4478_o;
  wire n4479_o;
  wire n4480_o;
  wire n4481_o;
  wire n4482_o;
  wire n4483_o;
  wire n4484_o;
  wire n4485_o;
  wire n4486_o;
  wire n4487_o;
  wire n4488_o;
  wire n4489_o;
  wire n4490_o;
  wire n4491_o;
  wire n4492_o;
  wire n4493_o;
  wire n4494_o;
  wire n4495_o;
  wire n4496_o;
  wire n4497_o;
  wire n4498_o;
  wire n4499_o;
  wire n4500_o;
  wire n4501_o;
  wire n4504_o;
  wire n4505_o;
  wire n4506_o;
  wire n4507_o;
  wire n4509_o;
  wire n4511_o;
  wire n4512_o;
  wire n4513_o;
  wire n4514_o;
  wire n4515_o;
  wire n4516_o;
  wire n4517_o;
  wire n4518_o;
  wire n4519_o;
  wire n4520_o;
  wire n4521_o;
  wire n4522_o;
  wire n4523_o;
  wire n4524_o;
  wire n4525_o;
  wire n4526_o;
  wire n4527_o;
  wire n4528_o;
  wire n4529_o;
  wire n4530_o;
  wire n4531_o;
  wire n4532_o;
  wire n4533_o;
  wire n4534_o;
  wire n4535_o;
  wire n4536_o;
  wire n4537_o;
  wire n4538_o;
  wire n4539_o;
  wire n4540_o;
  wire n4541_o;
  wire n4542_o;
  wire n4543_o;
  wire n4544_o;
  wire n4545_o;
  wire n4546_o;
  wire n4547_o;
  wire n4548_o;
  wire n4549_o;
  wire n4550_o;
  wire n4551_o;
  wire n4552_o;
  wire n4553_o;
  wire n4554_o;
  wire n4555_o;
  wire n4556_o;
  wire n4557_o;
  wire n4558_o;
  wire n4559_o;
  wire n4560_o;
  wire n4561_o;
  wire n4562_o;
  wire n4563_o;
  wire n4564_o;
  wire n4565_o;
  wire n4566_o;
  wire n4567_o;
  wire n4568_o;
  wire n4569_o;
  wire n4570_o;
  wire n4571_o;
  wire n4572_o;
  wire n4573_o;
  wire n4574_o;
  wire n4575_o;
  wire n4576_o;
  wire n4577_o;
  wire n4578_o;
  wire n4579_o;
  wire n4580_o;
  wire n4581_o;
  wire n4582_o;
  wire n4583_o;
  wire n4584_o;
  wire n4585_o;
  wire n4587_o;
  wire n4588_o;
  wire n4589_o;
  wire n4590_o;
  wire n4592_o;
  wire n4594_o;
  wire n4595_o;
  wire n4596_o;
  wire n4597_o;
  wire n4598_o;
  wire n4599_o;
  wire n4600_o;
  wire n4601_o;
  wire n4602_o;
  wire n4603_o;
  wire n4604_o;
  wire n4605_o;
  wire n4606_o;
  wire n4607_o;
  wire n4608_o;
  wire n4609_o;
  wire n4610_o;
  wire n4611_o;
  wire n4612_o;
  wire n4613_o;
  wire n4614_o;
  wire n4615_o;
  wire n4616_o;
  wire n4617_o;
  wire n4618_o;
  wire n4619_o;
  wire n4620_o;
  wire n4621_o;
  wire n4622_o;
  wire n4623_o;
  wire n4624_o;
  wire n4625_o;
  wire n4626_o;
  wire n4627_o;
  wire n4628_o;
  wire n4630_o;
  wire n4631_o;
  wire n4632_o;
  wire n4633_o;
  wire n4635_o;
  wire n4637_o;
  wire n4638_o;
  wire n4639_o;
  wire n4640_o;
  wire n4641_o;
  wire n4642_o;
  wire n4643_o;
  wire n4644_o;
  wire n4645_o;
  wire n4646_o;
  wire n4647_o;
  wire n4648_o;
  wire n4649_o;
  wire n4650_o;
  wire n4651_o;
  wire n4653_o;
  wire n4654_o;
  wire n4655_o;
  wire n4656_o;
  wire n4658_o;
  wire n4660_o;
  wire n4661_o;
  wire n4662_o;
  wire n4663_o;
  wire n4664_o;
  wire n4666_o;
  wire n4667_o;
  wire n4668_o;
  wire n4669_o;
  wire n4671_o;
  wire [5:0] n4673_o;
  wire [63:0] n4676_o;
  wire n4685_o;
  wire n4686_o;
  wire n4688_o;
  wire n4690_o;
  wire n4691_o;
  wire n4692_o;
  wire n4693_o;
  wire n4694_o;
  wire n4695_o;
  wire n4696_o;
  wire n4697_o;
  wire n4698_o;
  wire n4699_o;
  wire n4700_o;
  wire n4701_o;
  wire n4702_o;
  wire n4703_o;
  wire n4704_o;
  wire n4705_o;
  wire n4706_o;
  wire n4707_o;
  wire n4708_o;
  wire n4709_o;
  wire n4710_o;
  wire n4711_o;
  wire n4712_o;
  wire n4713_o;
  wire n4714_o;
  wire n4715_o;
  wire n4716_o;
  wire n4717_o;
  wire n4718_o;
  wire n4719_o;
  wire n4720_o;
  wire n4721_o;
  wire n4722_o;
  wire n4723_o;
  wire n4724_o;
  wire n4725_o;
  wire n4726_o;
  wire n4727_o;
  wire n4728_o;
  wire n4729_o;
  wire n4730_o;
  wire n4731_o;
  wire n4732_o;
  wire n4733_o;
  wire n4734_o;
  wire n4735_o;
  wire n4736_o;
  wire n4737_o;
  wire n4738_o;
  wire n4739_o;
  wire n4740_o;
  wire n4741_o;
  wire n4742_o;
  wire n4743_o;
  wire n4744_o;
  wire n4745_o;
  wire n4746_o;
  wire n4747_o;
  wire n4748_o;
  wire n4749_o;
  wire n4750_o;
  wire n4751_o;
  wire n4752_o;
  wire n4753_o;
  wire n4754_o;
  wire n4755_o;
  wire n4756_o;
  wire n4757_o;
  wire n4758_o;
  wire n4759_o;
  wire n4760_o;
  wire n4761_o;
  wire n4762_o;
  wire n4763_o;
  wire n4764_o;
  wire n4765_o;
  wire n4766_o;
  wire n4767_o;
  wire n4768_o;
  wire n4769_o;
  wire n4770_o;
  wire n4771_o;
  wire n4772_o;
  wire n4773_o;
  wire n4774_o;
  wire n4775_o;
  wire n4776_o;
  wire n4777_o;
  wire n4778_o;
  wire n4779_o;
  wire n4780_o;
  wire n4781_o;
  wire n4782_o;
  wire [1:0] n4785_o;
  wire n4786_o;
  wire n4788_o;
  wire [1:0] n4790_o;
  wire n4791_o;
  wire n4792_o;
  wire [1:0] n4793_o;
  wire n4794_o;
  wire n4795_o;
  wire [1:0] n4796_o;
  wire n4797_o;
  wire n4798_o;
  wire [1:0] n4799_o;
  wire n4800_o;
  wire n4801_o;
  wire [1:0] n4802_o;
  wire n4803_o;
  wire n4804_o;
  wire [1:0] n4805_o;
  wire n4806_o;
  wire n4807_o;
  wire [1:0] n4808_o;
  wire n4809_o;
  wire n4810_o;
  wire [1:0] n4811_o;
  wire n4812_o;
  wire n4813_o;
  wire [1:0] n4814_o;
  wire n4815_o;
  wire n4816_o;
  wire [1:0] n4817_o;
  wire n4818_o;
  wire n4819_o;
  wire [1:0] n4820_o;
  wire n4821_o;
  wire n4822_o;
  wire [1:0] n4823_o;
  wire n4824_o;
  wire n4825_o;
  wire [1:0] n4826_o;
  wire n4827_o;
  wire n4828_o;
  wire [1:0] n4829_o;
  wire n4830_o;
  wire n4831_o;
  wire [1:0] n4832_o;
  wire n4833_o;
  wire n4834_o;
  wire [3:0] n4836_o;
  wire n4837_o;
  wire n4839_o;
  wire [3:0] n4841_o;
  wire n4842_o;
  wire n4843_o;
  wire [3:0] n4844_o;
  wire n4845_o;
  wire n4846_o;
  wire [3:0] n4847_o;
  wire n4848_o;
  wire n4849_o;
  wire [3:0] n4850_o;
  wire n4851_o;
  wire n4852_o;
  wire [3:0] n4853_o;
  wire n4854_o;
  wire n4855_o;
  wire [3:0] n4856_o;
  wire n4857_o;
  wire n4858_o;
  wire [3:0] n4859_o;
  wire n4860_o;
  wire n4861_o;
  wire [7:0] n4863_o;
  wire n4864_o;
  wire n4866_o;
  wire [7:0] n4868_o;
  wire n4869_o;
  wire n4870_o;
  wire [7:0] n4871_o;
  wire n4872_o;
  wire n4873_o;
  wire [7:0] n4874_o;
  wire n4875_o;
  wire n4876_o;
  wire [15:0] n4878_o;
  wire n4879_o;
  wire n4881_o;
  wire [15:0] n4883_o;
  wire n4884_o;
  wire n4885_o;
  wire [31:0] n4887_o;
  wire n4888_o;
  wire n4890_o;
  wire [5:0] n4892_o;
  wire [3:0] n4894_o;
  wire [1:0] n4895_o;
  wire [5:0] n4896_o;
  wire [3:0] n4899_o;
  wire n4909_o;
  localparam [7:0] n4910_o = 8'b00000000;
  wire [4:0] n4911_o;
  wire [7:0] n4912_o;
  wire [7:0] n4914_o;
  reg [47:0] n4918_q;
  wire [11:0] n4919_o;
  reg [15:0] n4920_q;
  reg [32:0] n4921_q;
  wire [33:0] n4922_o;
  reg [11:0] n4923_q;
  wire n4924_o;
  wire n4925_o;
  wire n4926_o;
  wire n4927_o;
  wire n4928_o;
  wire n4929_o;
  wire n4930_o;
  wire n4931_o;
  wire n4932_o;
  wire n4933_o;
  wire n4934_o;
  wire n4935_o;
  wire n4936_o;
  wire n4937_o;
  wire n4938_o;
  wire n4939_o;
  wire [1:0] n4940_o;
  reg n4941_o;
  wire [1:0] n4942_o;
  reg n4943_o;
  wire [1:0] n4944_o;
  reg n4945_o;
  wire [1:0] n4946_o;
  reg n4947_o;
  wire [1:0] n4948_o;
  reg n4949_o;
  wire n4950_o;
  wire n4951_o;
  wire n4952_o;
  wire n4953_o;
  wire n4954_o;
  wire n4955_o;
  wire n4956_o;
  wire n4957_o;
  wire n4958_o;
  wire n4959_o;
  wire n4960_o;
  wire n4961_o;
  wire n4962_o;
  wire n4963_o;
  wire n4964_o;
  wire n4965_o;
  wire [1:0] n4966_o;
  reg n4967_o;
  wire [1:0] n4968_o;
  reg n4969_o;
  wire [1:0] n4970_o;
  reg n4971_o;
  wire [1:0] n4972_o;
  reg n4973_o;
  wire [1:0] n4974_o;
  reg n4975_o;
  wire [2:0] n4976_o;
  wire [2:0] n4977_o;
  wire [2:0] n4978_o;
  wire [2:0] n4979_o;
  wire [2:0] n4980_o;
  wire [2:0] n4981_o;
  wire [2:0] n4982_o;
  wire [2:0] n4983_o;
  wire [2:0] n4984_o;
  wire [2:0] n4985_o;
  wire [2:0] n4986_o;
  wire [2:0] n4987_o;
  wire [2:0] n4988_o;
  wire [2:0] n4989_o;
  wire [2:0] n4990_o;
  wire [2:0] n4991_o;
  wire [1:0] n4992_o;
  reg [2:0] n4993_o;
  wire [1:0] n4994_o;
  reg [2:0] n4995_o;
  wire [1:0] n4996_o;
  reg [2:0] n4997_o;
  wire [1:0] n4998_o;
  reg [2:0] n4999_o;
  wire [1:0] n5000_o;
  reg [2:0] n5001_o;
  wire n5002_o;
  wire n5003_o;
  wire n5004_o;
  wire n5005_o;
  wire n5006_o;
  wire n5007_o;
  wire n5008_o;
  wire n5009_o;
  wire n5010_o;
  wire n5011_o;
  wire n5012_o;
  wire n5013_o;
  wire n5014_o;
  wire n5015_o;
  wire n5016_o;
  wire n5017_o;
  wire n5018_o;
  wire n5019_o;
  wire n5020_o;
  wire n5021_o;
  wire n5022_o;
  wire n5023_o;
  wire n5024_o;
  wire n5025_o;
  wire n5026_o;
  wire n5027_o;
  wire n5028_o;
  wire n5029_o;
  wire n5030_o;
  wire n5031_o;
  wire n5032_o;
  wire n5033_o;
  wire n5034_o;
  wire n5035_o;
  wire n5036_o;
  wire n5037_o;
  wire [2:0] n5038_o;
  wire [2:0] n5039_o;
  wire [2:0] n5040_o;
  wire [2:0] n5041_o;
  wire [2:0] n5042_o;
  wire [2:0] n5043_o;
  wire [2:0] n5044_o;
  wire [2:0] n5045_o;
  wire [2:0] n5046_o;
  wire [2:0] n5047_o;
  wire [2:0] n5048_o;
  wire [2:0] n5049_o;
  wire [2:0] n5050_o;
  wire [2:0] n5051_o;
  wire [2:0] n5052_o;
  wire [2:0] n5053_o;
  wire [2:0] n5054_o;
  wire [2:0] n5055_o;
  wire [2:0] n5056_o;
  wire [2:0] n5057_o;
  wire [2:0] n5058_o;
  wire [2:0] n5059_o;
  wire [2:0] n5060_o;
  wire [2:0] n5061_o;
  wire [2:0] n5062_o;
  wire [2:0] n5063_o;
  wire [2:0] n5064_o;
  wire [2:0] n5065_o;
  wire [2:0] n5066_o;
  wire [2:0] n5067_o;
  wire [2:0] n5068_o;
  wire [2:0] n5069_o;
  wire [47:0] n5070_o;
  wire n5071_o;
  wire n5072_o;
  wire n5073_o;
  wire n5074_o;
  wire n5075_o;
  wire n5076_o;
  wire n5077_o;
  wire n5078_o;
  wire n5079_o;
  wire n5080_o;
  wire n5081_o;
  wire n5082_o;
  wire n5083_o;
  wire n5084_o;
  wire n5085_o;
  wire n5086_o;
  wire n5087_o;
  wire n5088_o;
  wire n5089_o;
  wire n5090_o;
  wire n5091_o;
  wire n5092_o;
  wire n5093_o;
  wire n5094_o;
  wire n5095_o;
  wire n5096_o;
  wire n5097_o;
  wire n5098_o;
  wire n5099_o;
  wire n5100_o;
  wire n5101_o;
  wire n5102_o;
  wire n5103_o;
  wire n5104_o;
  wire [7:0] n5105_o;
  wire n5106_o;
  wire n5107_o;
  wire n5108_o;
  wire n5109_o;
  wire n5110_o;
  wire n5111_o;
  wire n5112_o;
  wire n5113_o;
  wire n5114_o;
  wire n5115_o;
  wire n5116_o;
  wire n5117_o;
  wire n5118_o;
  wire n5119_o;
  wire n5120_o;
  wire n5121_o;
  wire n5122_o;
  wire n5123_o;
  wire n5124_o;
  wire n5125_o;
  wire n5126_o;
  wire n5127_o;
  wire n5128_o;
  wire n5129_o;
  wire n5130_o;
  wire n5131_o;
  wire n5132_o;
  wire n5133_o;
  wire n5134_o;
  wire n5135_o;
  wire n5136_o;
  wire n5137_o;
  wire n5138_o;
  wire n5139_o;
  wire [7:0] n5140_o;
  wire n5141_o;
  wire n5142_o;
  wire n5143_o;
  wire n5144_o;
  wire n5145_o;
  wire n5146_o;
  wire n5147_o;
  wire n5148_o;
  wire n5149_o;
  wire n5150_o;
  wire n5151_o;
  wire n5152_o;
  wire n5153_o;
  wire n5154_o;
  wire n5155_o;
  wire n5156_o;
  wire n5157_o;
  wire n5158_o;
  wire n5159_o;
  wire n5160_o;
  wire n5161_o;
  wire n5162_o;
  wire n5163_o;
  wire n5164_o;
  wire n5165_o;
  wire n5166_o;
  wire n5167_o;
  wire n5168_o;
  wire n5169_o;
  wire n5170_o;
  wire n5171_o;
  wire n5172_o;
  wire n5173_o;
  wire n5174_o;
  wire [7:0] n5175_o;
  wire n5176_o;
  wire n5177_o;
  wire n5178_o;
  wire n5179_o;
  wire n5180_o;
  wire n5181_o;
  wire n5182_o;
  wire n5183_o;
  wire n5184_o;
  wire n5185_o;
  wire n5186_o;
  wire n5187_o;
  wire n5188_o;
  wire n5189_o;
  wire n5190_o;
  wire n5191_o;
  wire n5192_o;
  wire n5193_o;
  wire n5194_o;
  wire n5195_o;
  wire n5196_o;
  wire n5197_o;
  wire n5198_o;
  wire n5199_o;
  wire n5200_o;
  wire n5201_o;
  wire n5202_o;
  wire n5203_o;
  wire n5204_o;
  wire n5205_o;
  wire n5206_o;
  wire n5207_o;
  wire n5208_o;
  wire n5209_o;
  wire [7:0] n5210_o;
  wire n5211_o;
  wire n5212_o;
  wire n5213_o;
  wire n5214_o;
  wire n5215_o;
  wire n5216_o;
  wire n5217_o;
  wire n5218_o;
  wire n5219_o;
  wire n5220_o;
  wire n5221_o;
  wire n5222_o;
  wire n5223_o;
  wire n5224_o;
  wire n5225_o;
  wire n5226_o;
  wire n5227_o;
  wire n5228_o;
  wire n5229_o;
  wire n5230_o;
  wire n5231_o;
  wire n5232_o;
  wire n5233_o;
  wire n5234_o;
  wire n5235_o;
  wire n5236_o;
  wire n5237_o;
  wire n5238_o;
  wire n5239_o;
  wire n5240_o;
  wire n5241_o;
  wire n5242_o;
  wire n5243_o;
  wire n5244_o;
  wire [7:0] n5245_o;
  wire n5246_o;
  wire n5247_o;
  wire n5248_o;
  wire n5249_o;
  wire n5250_o;
  wire n5251_o;
  wire n5252_o;
  wire n5253_o;
  wire n5254_o;
  wire n5255_o;
  wire n5256_o;
  wire n5257_o;
  wire n5258_o;
  wire n5259_o;
  wire n5260_o;
  wire n5261_o;
  wire n5262_o;
  wire n5263_o;
  wire n5264_o;
  wire n5265_o;
  wire n5266_o;
  wire n5267_o;
  wire n5268_o;
  wire n5269_o;
  wire n5270_o;
  wire n5271_o;
  wire n5272_o;
  wire n5273_o;
  wire n5274_o;
  wire n5275_o;
  wire n5276_o;
  wire n5277_o;
  wire n5278_o;
  wire n5279_o;
  wire [7:0] n5280_o;
  wire n5281_o;
  wire n5282_o;
  wire n5283_o;
  wire n5284_o;
  wire n5285_o;
  wire n5286_o;
  wire n5287_o;
  wire n5288_o;
  wire n5289_o;
  wire n5290_o;
  wire n5291_o;
  wire n5292_o;
  wire n5293_o;
  wire n5294_o;
  wire n5295_o;
  wire n5296_o;
  wire n5297_o;
  wire n5298_o;
  wire n5299_o;
  wire n5300_o;
  wire n5301_o;
  wire n5302_o;
  wire n5303_o;
  wire n5304_o;
  wire n5305_o;
  wire n5306_o;
  wire n5307_o;
  wire n5308_o;
  wire n5309_o;
  wire n5310_o;
  wire n5311_o;
  wire n5312_o;
  wire n5313_o;
  wire n5314_o;
  wire [7:0] n5315_o;
  wire n5316_o;
  wire n5317_o;
  wire n5318_o;
  wire n5319_o;
  wire n5320_o;
  wire n5321_o;
  wire n5322_o;
  wire n5323_o;
  wire n5324_o;
  wire n5325_o;
  wire n5326_o;
  wire n5327_o;
  wire n5328_o;
  wire n5329_o;
  wire n5330_o;
  wire n5331_o;
  wire n5332_o;
  wire n5333_o;
  wire n5334_o;
  wire n5335_o;
  wire n5336_o;
  wire n5337_o;
  wire n5338_o;
  wire n5339_o;
  wire n5340_o;
  wire n5341_o;
  wire n5342_o;
  wire n5343_o;
  wire n5344_o;
  wire n5345_o;
  wire n5346_o;
  wire n5347_o;
  wire n5348_o;
  wire n5349_o;
  wire [7:0] n5350_o;
  wire n5351_o;
  wire n5352_o;
  wire n5353_o;
  wire n5354_o;
  wire n5355_o;
  wire n5356_o;
  wire n5357_o;
  wire n5358_o;
  wire n5359_o;
  wire n5360_o;
  wire n5361_o;
  wire n5362_o;
  wire n5363_o;
  wire n5364_o;
  wire n5365_o;
  wire n5366_o;
  wire n5367_o;
  wire n5368_o;
  wire n5369_o;
  wire n5370_o;
  wire n5371_o;
  wire n5372_o;
  wire n5373_o;
  wire n5374_o;
  wire n5375_o;
  wire n5376_o;
  wire n5377_o;
  wire n5378_o;
  wire n5379_o;
  wire n5380_o;
  wire n5381_o;
  wire n5382_o;
  wire n5383_o;
  wire n5384_o;
  wire [7:0] n5385_o;
  wire n5386_o;
  wire n5387_o;
  wire n5388_o;
  wire n5389_o;
  wire n5390_o;
  wire n5391_o;
  wire n5392_o;
  wire n5393_o;
  wire n5394_o;
  wire n5395_o;
  wire n5396_o;
  wire n5397_o;
  wire n5398_o;
  wire n5399_o;
  wire n5400_o;
  wire n5401_o;
  wire n5402_o;
  wire n5403_o;
  wire n5404_o;
  wire n5405_o;
  wire n5406_o;
  wire n5407_o;
  wire n5408_o;
  wire n5409_o;
  wire n5410_o;
  wire n5411_o;
  wire n5412_o;
  wire n5413_o;
  wire n5414_o;
  wire n5415_o;
  wire n5416_o;
  wire n5417_o;
  wire n5418_o;
  wire n5419_o;
  wire [7:0] n5420_o;
  wire n5421_o;
  wire n5422_o;
  wire n5423_o;
  wire n5424_o;
  wire n5425_o;
  wire n5426_o;
  wire n5427_o;
  wire n5428_o;
  wire n5429_o;
  wire n5430_o;
  wire n5431_o;
  wire n5432_o;
  wire n5433_o;
  wire n5434_o;
  wire n5435_o;
  wire n5436_o;
  wire n5437_o;
  wire n5438_o;
  wire n5439_o;
  wire n5440_o;
  wire n5441_o;
  wire n5442_o;
  wire n5443_o;
  wire n5444_o;
  wire n5445_o;
  wire n5446_o;
  wire n5447_o;
  wire n5448_o;
  wire n5449_o;
  wire n5450_o;
  wire n5451_o;
  wire n5452_o;
  wire n5453_o;
  wire n5454_o;
  wire [7:0] n5455_o;
  wire n5456_o;
  wire n5457_o;
  wire n5458_o;
  wire n5459_o;
  wire n5460_o;
  wire n5461_o;
  wire n5462_o;
  wire n5463_o;
  wire n5464_o;
  wire n5465_o;
  wire n5466_o;
  wire n5467_o;
  wire n5468_o;
  wire n5469_o;
  wire n5470_o;
  wire n5471_o;
  wire n5472_o;
  wire n5473_o;
  wire n5474_o;
  wire n5475_o;
  wire n5476_o;
  wire n5477_o;
  wire n5478_o;
  wire n5479_o;
  wire n5480_o;
  wire n5481_o;
  wire n5482_o;
  wire n5483_o;
  wire n5484_o;
  wire n5485_o;
  wire n5486_o;
  wire n5487_o;
  wire n5488_o;
  wire n5489_o;
  wire [7:0] n5490_o;
  wire n5491_o;
  wire n5492_o;
  wire n5493_o;
  wire n5494_o;
  wire n5495_o;
  wire n5496_o;
  wire n5497_o;
  wire n5498_o;
  wire n5499_o;
  wire n5500_o;
  wire n5501_o;
  wire n5502_o;
  wire n5503_o;
  wire n5504_o;
  wire n5505_o;
  wire n5506_o;
  wire n5507_o;
  wire n5508_o;
  wire n5509_o;
  wire n5510_o;
  wire n5511_o;
  wire n5512_o;
  wire n5513_o;
  wire n5514_o;
  wire n5515_o;
  wire n5516_o;
  wire n5517_o;
  wire n5518_o;
  wire n5519_o;
  wire n5520_o;
  wire n5521_o;
  wire n5522_o;
  wire n5523_o;
  wire n5524_o;
  wire [7:0] n5525_o;
  wire n5526_o;
  wire n5527_o;
  wire n5528_o;
  wire n5529_o;
  wire n5530_o;
  wire n5531_o;
  wire n5532_o;
  wire n5533_o;
  wire n5534_o;
  wire n5535_o;
  wire n5536_o;
  wire n5537_o;
  wire n5538_o;
  wire n5539_o;
  wire n5540_o;
  wire n5541_o;
  wire n5542_o;
  wire n5543_o;
  wire n5544_o;
  wire n5545_o;
  wire n5546_o;
  wire n5547_o;
  wire n5548_o;
  wire n5549_o;
  wire n5550_o;
  wire n5551_o;
  wire n5552_o;
  wire n5553_o;
  wire n5554_o;
  wire n5555_o;
  wire n5556_o;
  wire n5557_o;
  wire n5558_o;
  wire n5559_o;
  wire [7:0] n5560_o;
  wire n5561_o;
  wire n5562_o;
  wire n5563_o;
  wire n5564_o;
  wire n5565_o;
  wire n5566_o;
  wire n5567_o;
  wire n5568_o;
  wire n5569_o;
  wire n5570_o;
  wire n5571_o;
  wire n5572_o;
  wire n5573_o;
  wire n5574_o;
  wire n5575_o;
  wire n5576_o;
  wire n5577_o;
  wire n5578_o;
  wire n5579_o;
  wire n5580_o;
  wire n5581_o;
  wire n5582_o;
  wire n5583_o;
  wire n5584_o;
  wire n5585_o;
  wire n5586_o;
  wire n5587_o;
  wire n5588_o;
  wire n5589_o;
  wire n5590_o;
  wire n5591_o;
  wire n5592_o;
  wire n5593_o;
  wire n5594_o;
  wire [7:0] n5595_o;
  wire n5596_o;
  wire n5597_o;
  wire n5598_o;
  wire n5599_o;
  wire n5600_o;
  wire n5601_o;
  wire n5602_o;
  wire n5603_o;
  wire n5604_o;
  wire n5605_o;
  wire n5606_o;
  wire n5607_o;
  wire n5608_o;
  wire n5609_o;
  wire n5610_o;
  wire n5611_o;
  wire n5612_o;
  wire n5613_o;
  wire n5614_o;
  wire n5615_o;
  wire n5616_o;
  wire n5617_o;
  wire n5618_o;
  wire n5619_o;
  wire n5620_o;
  wire n5621_o;
  wire n5622_o;
  wire n5623_o;
  wire n5624_o;
  wire n5625_o;
  wire n5626_o;
  wire n5627_o;
  wire n5628_o;
  wire n5629_o;
  wire [7:0] n5630_o;
  assign wb_out_dat = n3083_o;
  assign wb_out_ack = n3084_o;
  assign wb_out_stall = n3085_o;
  assign icp_out_src = n3087_o;
  assign icp_out_pri = n3088_o;
  /* xics.vhdl:36:9  */
  assign n3081_o = {wb_in_we, wb_in_stb, wb_in_cyc, wb_in_sel, wb_in_dat, wb_in_adr};
  assign n3083_o = n4922_o[31:0];
  /* xics.vhdl:187:17  */
  assign n3084_o = n4922_o[32];
  /* xics.vhdl:183:22  */
  assign n3085_o = n4922_o[33];
  assign n3087_o = n4923_q[3:0];
  assign n3088_o = n4923_q[11:4];
  /* xics.vhdl:241:12  */
  assign xives = n4918_q; // (signal)
  /* xics.vhdl:243:12  */
  assign wb_valid = n3111_o; // (signal)
  /* xics.vhdl:244:12  */
  assign reg_idx = n3102_o; // (signal)
  /* xics.vhdl:245:12  */
  assign icp_out_next = n4919_o; // (signal)
  /* xics.vhdl:246:12  */
  assign int_level_l = n4920_q; // (signal)
  /* xics.vhdl:332:12  */
  assign reg_is_xive = n3089_o; // (signal)
  /* xics.vhdl:333:12  */
  assign reg_is_config = n3094_o; // (signal)
  /* xics.vhdl:334:12  */
  assign reg_is_debug = n3100_o; // (signal)
  /* xics.vhdl:340:31  */
  assign n3089_o = n3081_o[9];
  /* xics.vhdl:341:40  */
  assign n3091_o = n3081_o[9:0];
  /* xics.vhdl:341:53  */
  assign n3093_o = n3091_o == 10'b0000000000;
  /* xics.vhdl:341:26  */
  assign n3094_o = n3093_o ? 1'b1 : 1'b0;
  /* xics.vhdl:342:40  */
  assign n3097_o = n3081_o[9:0];
  /* xics.vhdl:342:53  */
  assign n3099_o = n3097_o == 10'b0000000001;
  /* xics.vhdl:342:26  */
  assign n3100_o = n3099_o ? 1'b1 : 1'b0;
  /* xics.vhdl:345:45  */
  assign n3102_o = n3081_o[3:0];
  /* xics.vhdl:358:23  */
  assign n3109_o = n3081_o[66];
  /* xics.vhdl:358:37  */
  assign n3110_o = n3081_o[67];
  /* xics.vhdl:358:27  */
  assign n3111_o = n3109_o & n3110_o;
  /* xics.vhdl:369:48  */
  assign n3118_o = {n4949_o, 1'b0};
  /* xics.vhdl:370:31  */
  assign n3121_o = {n3118_o, n4975_o};
  /* xics.vhdl:371:48  */
  assign n3123_o = {n3121_o, 1'b0};
  /* xics.vhdl:372:31  */
  assign n3125_o = {n3123_o, 20'b00000000000000000000};
  /* xics.vhdl:374:45  */
  assign n3128_o = 4'b1111 - reg_idx;
  /* xics.vhdl:374:54  */
  assign n3131_o = n5001_o[2:0];
  /* xics.vhdl:282:16  */
  assign n3138_o = n3131_o == 3'b111;
  assign n3140_o = n3139_o[7:3];
  assign n3141_o = {n3140_o, n3131_o};
  /* xics.vhdl:282:9  */
  assign n3143_o = n3138_o ? 8'b11111111 : n3141_o;
  /* xics.vhdl:373:36  */
  assign n3145_o = {n3125_o, n3143_o};
  /* xics.vhdl:378:51  */
  assign n3147_o = icp_out_next[3:0];
  /* xics.vhdl:378:36  */
  assign n3149_o = {20'b00000000000000000000, n3147_o};
  /* xics.vhdl:378:70  */
  assign n3150_o = icp_out_next[11:4];
  /* xics.vhdl:378:55  */
  assign n3151_o = {n3149_o, n3150_o};
  /* xics.vhdl:377:13  */
  assign n3153_o = reg_is_debug ? n3151_o : 32'b00000000000000000000000000000000;
  /* xics.vhdl:375:13  */
  assign n3155_o = reg_is_config ? 32'b00000011000000000000000000010000 : n3153_o;
  /* xics.vhdl:368:13  */
  assign n3156_o = reg_is_xive ? n3145_o : n3155_o;
  /* xics.vhdl:251:29  */
  assign n3164_o = n3156_o[31:24];
  /* xics.vhdl:252:29  */
  assign n3167_o = n3156_o[23:16];
  /* xics.vhdl:253:29  */
  assign n3169_o = n3156_o[15:8];
  /* xics.vhdl:254:29  */
  assign n3171_o = n3156_o[7:0];
  assign n3172_o = {n3171_o, n3169_o, n3167_o, n3164_o};
  assign n3173_o = {wb_valid, n3172_o};
  /* xics.vhdl:390:30  */
  assign n3181_o = n3081_o[61:30];
  /* xics.vhdl:251:29  */
  assign n3187_o = n3181_o[31:24];
  /* xics.vhdl:252:29  */
  assign n3190_o = n3181_o[23:16];
  /* xics.vhdl:253:29  */
  assign n3192_o = n3181_o[15:8];
  /* xics.vhdl:254:29  */
  assign n3194_o = n3181_o[7:0];
  assign n3195_o = {n3194_o, n3192_o, n3190_o, n3187_o};
  /* xics.vhdl:397:44  */
  assign n3213_o = n3081_o[68];
  /* xics.vhdl:397:34  */
  assign n3214_o = wb_valid & n3213_o;
  /* xics.vhdl:401:27  */
  assign n3216_o = 4'b1111 - reg_idx;
  /* xics.vhdl:401:58  */
  assign n3219_o = n3195_o[7:0];
  assign n3227_o = n3226_o[7:3];
  assign n3228_o = {n3227_o, 3'b111};
  /* xics.vhdl:272:27  */
  assign n3229_o = $unsigned(n3219_o) >= $unsigned(n3228_o);
  /* xics.vhdl:275:24  */
  assign n3231_o = n3219_o[2:0];
  /* xics.vhdl:272:9  */
  assign n3232_o = n3229_o ? 3'b111 : n3231_o;
  /* xics.vhdl:397:13  */
  assign n3234_o = n3235_o ? n5070_o : xives;
  /* xics.vhdl:397:13  */
  assign n3235_o = n3214_o & reg_is_xive;
  assign n3236_o = {3'b111, 3'b111, 3'b111, 3'b111, 3'b111, 3'b111, 3'b111, 3'b111, 3'b111, 3'b111, 3'b111, 3'b111, 3'b111, 3'b111, 3'b111, 3'b111};
  /* xics.vhdl:393:13  */
  assign n3237_o = rst ? n3236_o : n3234_o;
  /* xics.vhdl:431:27  */
  assign n3249_o = int_level_l[0];
  /* xics.vhdl:432:64  */
  assign n3251_o = xives[47:45];
  /* xics.vhdl:432:68  */
  assign n3252_o = n3251_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3265_o = 8'b00000000 | n5105_o;
  /* xics.vhdl:431:13  */
  assign n3267_o = n3249_o ? n3265_o : 8'b00000000;
  /* xics.vhdl:431:27  */
  assign n3269_o = int_level_l[1];
  /* xics.vhdl:432:64  */
  assign n3271_o = xives[44:42];
  /* xics.vhdl:432:68  */
  assign n3272_o = n3271_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3284_o = n3267_o | n5140_o;
  /* xics.vhdl:431:13  */
  assign n3285_o = n3269_o ? n3284_o : n3267_o;
  /* xics.vhdl:431:27  */
  assign n3286_o = int_level_l[2];
  /* xics.vhdl:432:64  */
  assign n3288_o = xives[41:39];
  /* xics.vhdl:432:68  */
  assign n3289_o = n3288_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3301_o = n3285_o | n5175_o;
  /* xics.vhdl:431:13  */
  assign n3302_o = n3286_o ? n3301_o : n3285_o;
  /* xics.vhdl:431:27  */
  assign n3303_o = int_level_l[3];
  /* xics.vhdl:432:64  */
  assign n3305_o = xives[38:36];
  /* xics.vhdl:432:68  */
  assign n3306_o = n3305_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3318_o = n3302_o | n5210_o;
  /* xics.vhdl:431:13  */
  assign n3319_o = n3303_o ? n3318_o : n3302_o;
  /* xics.vhdl:431:27  */
  assign n3320_o = int_level_l[4];
  /* xics.vhdl:432:64  */
  assign n3322_o = xives[35:33];
  /* xics.vhdl:432:68  */
  assign n3323_o = n3322_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3335_o = n3319_o | n5245_o;
  /* xics.vhdl:431:13  */
  assign n3336_o = n3320_o ? n3335_o : n3319_o;
  /* xics.vhdl:431:27  */
  assign n3337_o = int_level_l[5];
  /* xics.vhdl:432:64  */
  assign n3339_o = xives[32:30];
  /* xics.vhdl:432:68  */
  assign n3340_o = n3339_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3352_o = n3336_o | n5280_o;
  /* xics.vhdl:431:13  */
  assign n3353_o = n3337_o ? n3352_o : n3336_o;
  /* xics.vhdl:431:27  */
  assign n3354_o = int_level_l[6];
  /* xics.vhdl:432:64  */
  assign n3356_o = xives[29:27];
  /* xics.vhdl:432:68  */
  assign n3357_o = n3356_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3369_o = n3353_o | n5315_o;
  /* xics.vhdl:431:13  */
  assign n3370_o = n3354_o ? n3369_o : n3353_o;
  /* xics.vhdl:431:27  */
  assign n3371_o = int_level_l[7];
  /* xics.vhdl:432:64  */
  assign n3373_o = xives[26:24];
  /* xics.vhdl:432:68  */
  assign n3374_o = n3373_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3386_o = n3370_o | n5350_o;
  /* xics.vhdl:431:13  */
  assign n3387_o = n3371_o ? n3386_o : n3370_o;
  /* xics.vhdl:431:27  */
  assign n3388_o = int_level_l[8];
  /* xics.vhdl:432:64  */
  assign n3390_o = xives[23:21];
  /* xics.vhdl:432:68  */
  assign n3391_o = n3390_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3403_o = n3387_o | n5385_o;
  /* xics.vhdl:431:13  */
  assign n3404_o = n3388_o ? n3403_o : n3387_o;
  /* xics.vhdl:431:27  */
  assign n3405_o = int_level_l[9];
  /* xics.vhdl:432:64  */
  assign n3407_o = xives[20:18];
  /* xics.vhdl:432:68  */
  assign n3408_o = n3407_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3420_o = n3404_o | n5420_o;
  /* xics.vhdl:431:13  */
  assign n3421_o = n3405_o ? n3420_o : n3404_o;
  /* xics.vhdl:431:27  */
  assign n3422_o = int_level_l[10];
  /* xics.vhdl:432:64  */
  assign n3424_o = xives[17:15];
  /* xics.vhdl:432:68  */
  assign n3425_o = n3424_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3437_o = n3421_o | n5455_o;
  /* xics.vhdl:431:13  */
  assign n3438_o = n3422_o ? n3437_o : n3421_o;
  /* xics.vhdl:431:27  */
  assign n3439_o = int_level_l[11];
  /* xics.vhdl:432:64  */
  assign n3441_o = xives[14:12];
  /* xics.vhdl:432:68  */
  assign n3442_o = n3441_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3454_o = n3438_o | n5490_o;
  /* xics.vhdl:431:13  */
  assign n3455_o = n3439_o ? n3454_o : n3438_o;
  /* xics.vhdl:431:27  */
  assign n3456_o = int_level_l[12];
  /* xics.vhdl:432:64  */
  assign n3458_o = xives[11:9];
  /* xics.vhdl:432:68  */
  assign n3459_o = n3458_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3471_o = n3455_o | n5525_o;
  /* xics.vhdl:431:13  */
  assign n3472_o = n3456_o ? n3471_o : n3455_o;
  /* xics.vhdl:431:27  */
  assign n3473_o = int_level_l[13];
  /* xics.vhdl:432:64  */
  assign n3475_o = xives[8:6];
  /* xics.vhdl:432:68  */
  assign n3476_o = n3475_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3488_o = n3472_o | n5560_o;
  /* xics.vhdl:431:13  */
  assign n3489_o = n3473_o ? n3488_o : n3472_o;
  /* xics.vhdl:431:27  */
  assign n3490_o = int_level_l[14];
  /* xics.vhdl:432:64  */
  assign n3492_o = xives[5:3];
  /* xics.vhdl:432:68  */
  assign n3493_o = n3492_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3505_o = n3489_o | n5595_o;
  /* xics.vhdl:431:13  */
  assign n3506_o = n3490_o ? n3505_o : n3489_o;
  /* xics.vhdl:431:27  */
  assign n3507_o = int_level_l[15];
  /* xics.vhdl:432:64  */
  assign n3509_o = xives[2:0];
  /* xics.vhdl:432:68  */
  assign n3510_o = n3509_o[2:0];
  /* xics.vhdl:432:44  */
  assign n3522_o = n3506_o | n5630_o;
  assign n3533_o = n3522_o[6:0];
  assign n3534_o = n3505_o[6:0];
  assign n3535_o = n3488_o[6:0];
  assign n3536_o = n3471_o[6:0];
  assign n3537_o = n3454_o[6:0];
  assign n3538_o = n3437_o[6:0];
  assign n3539_o = n3420_o[6:0];
  assign n3540_o = n3403_o[6:0];
  assign n3541_o = n3386_o[6:0];
  assign n3542_o = n3369_o[6:0];
  assign n3543_o = n3352_o[6:0];
  assign n3544_o = n3335_o[6:0];
  assign n3545_o = n3318_o[6:0];
  assign n3546_o = n3301_o[6:0];
  assign n3547_o = n3284_o[6:0];
  assign n3548_o = n3265_o[6:0];
  assign n3549_o = n3266_o[6:0];
  /* xics.vhdl:431:13  */
  assign n3550_o = n3249_o ? n3548_o : n3549_o;
  /* xics.vhdl:431:13  */
  assign n3551_o = n3269_o ? n3547_o : n3550_o;
  /* xics.vhdl:431:13  */
  assign n3552_o = n3286_o ? n3546_o : n3551_o;
  /* xics.vhdl:431:13  */
  assign n3553_o = n3303_o ? n3545_o : n3552_o;
  /* xics.vhdl:431:13  */
  assign n3554_o = n3320_o ? n3544_o : n3553_o;
  /* xics.vhdl:431:13  */
  assign n3555_o = n3337_o ? n3543_o : n3554_o;
  /* xics.vhdl:431:13  */
  assign n3556_o = n3354_o ? n3542_o : n3555_o;
  /* xics.vhdl:431:13  */
  assign n3557_o = n3371_o ? n3541_o : n3556_o;
  /* xics.vhdl:431:13  */
  assign n3558_o = n3388_o ? n3540_o : n3557_o;
  /* xics.vhdl:431:13  */
  assign n3559_o = n3405_o ? n3539_o : n3558_o;
  /* xics.vhdl:431:13  */
  assign n3560_o = n3422_o ? n3538_o : n3559_o;
  /* xics.vhdl:431:13  */
  assign n3561_o = n3439_o ? n3537_o : n3560_o;
  /* xics.vhdl:431:13  */
  assign n3562_o = n3456_o ? n3536_o : n3561_o;
  /* xics.vhdl:431:13  */
  assign n3563_o = n3473_o ? n3535_o : n3562_o;
  /* xics.vhdl:431:13  */
  assign n3564_o = n3490_o ? n3534_o : n3563_o;
  /* xics.vhdl:431:13  */
  assign n3565_o = n3507_o ? n3533_o : n3564_o;
  assign n3577_o = {1'b1, n3565_o};
  /* helpers.vhdl:282:34  */
  assign n3578_o = -n3577_o;
  assign n3580_o = {1'b1, n3565_o};
  /* helpers.vhdl:283:23  */
  assign n3581_o = n3578_o & n3580_o;
  assign n3583_o = {1'b1, n3565_o};
  /* helpers.vhdl:284:21  */
  assign n3584_o = n3578_o | n3583_o;
  /* helpers.vhdl:285:48  */
  assign n3587_o = {{56{n3584_o[7]}}, n3584_o}; // sext
  /* helpers.vhdl:266:29  */
  assign n3596_o = n3587_o[1];
  /* helpers.vhdl:266:55  */
  assign n3597_o = n3587_o[0];
  /* helpers.vhdl:266:50  */
  assign n3598_o = ~n3597_o;
  /* helpers.vhdl:266:46  */
  assign n3599_o = n3596_o & n3598_o;
  /* helpers.vhdl:266:24  */
  assign n3601_o = 1'b0 | n3599_o;
  /* helpers.vhdl:266:29  */
  assign n3603_o = n3587_o[3];
  /* helpers.vhdl:266:55  */
  assign n3604_o = n3587_o[2];
  /* helpers.vhdl:266:50  */
  assign n3605_o = ~n3604_o;
  /* helpers.vhdl:266:46  */
  assign n3606_o = n3603_o & n3605_o;
  /* helpers.vhdl:266:24  */
  assign n3607_o = n3601_o | n3606_o;
  /* helpers.vhdl:266:29  */
  assign n3608_o = n3587_o[5];
  /* helpers.vhdl:266:55  */
  assign n3609_o = n3587_o[4];
  /* helpers.vhdl:266:50  */
  assign n3610_o = ~n3609_o;
  /* helpers.vhdl:266:46  */
  assign n3611_o = n3608_o & n3610_o;
  /* helpers.vhdl:266:24  */
  assign n3612_o = n3607_o | n3611_o;
  /* helpers.vhdl:266:29  */
  assign n3613_o = n3587_o[7];
  /* helpers.vhdl:266:55  */
  assign n3614_o = n3587_o[6];
  /* helpers.vhdl:266:50  */
  assign n3615_o = ~n3614_o;
  /* helpers.vhdl:266:46  */
  assign n3616_o = n3613_o & n3615_o;
  /* helpers.vhdl:266:24  */
  assign n3617_o = n3612_o | n3616_o;
  /* helpers.vhdl:266:29  */
  assign n3618_o = n3587_o[9];
  /* helpers.vhdl:266:55  */
  assign n3619_o = n3587_o[8];
  /* helpers.vhdl:266:50  */
  assign n3620_o = ~n3619_o;
  /* helpers.vhdl:266:46  */
  assign n3621_o = n3618_o & n3620_o;
  /* helpers.vhdl:266:24  */
  assign n3622_o = n3617_o | n3621_o;
  /* helpers.vhdl:266:29  */
  assign n3623_o = n3587_o[11];
  /* helpers.vhdl:266:55  */
  assign n3624_o = n3587_o[10];
  /* helpers.vhdl:266:50  */
  assign n3625_o = ~n3624_o;
  /* helpers.vhdl:266:46  */
  assign n3626_o = n3623_o & n3625_o;
  /* helpers.vhdl:266:24  */
  assign n3627_o = n3622_o | n3626_o;
  /* helpers.vhdl:266:29  */
  assign n3628_o = n3587_o[13];
  /* helpers.vhdl:266:55  */
  assign n3629_o = n3587_o[12];
  /* helpers.vhdl:266:50  */
  assign n3630_o = ~n3629_o;
  /* helpers.vhdl:266:46  */
  assign n3631_o = n3628_o & n3630_o;
  /* helpers.vhdl:266:24  */
  assign n3632_o = n3627_o | n3631_o;
  /* helpers.vhdl:266:29  */
  assign n3633_o = n3587_o[15];
  /* helpers.vhdl:266:55  */
  assign n3634_o = n3587_o[14];
  /* helpers.vhdl:266:50  */
  assign n3635_o = ~n3634_o;
  /* helpers.vhdl:266:46  */
  assign n3636_o = n3633_o & n3635_o;
  /* helpers.vhdl:266:24  */
  assign n3637_o = n3632_o | n3636_o;
  /* helpers.vhdl:266:29  */
  assign n3638_o = n3587_o[17];
  /* helpers.vhdl:266:55  */
  assign n3639_o = n3587_o[16];
  /* helpers.vhdl:266:50  */
  assign n3640_o = ~n3639_o;
  /* helpers.vhdl:266:46  */
  assign n3641_o = n3638_o & n3640_o;
  /* helpers.vhdl:266:24  */
  assign n3642_o = n3637_o | n3641_o;
  /* helpers.vhdl:266:29  */
  assign n3643_o = n3587_o[19];
  /* helpers.vhdl:266:55  */
  assign n3644_o = n3587_o[18];
  /* helpers.vhdl:266:50  */
  assign n3645_o = ~n3644_o;
  /* helpers.vhdl:266:46  */
  assign n3646_o = n3643_o & n3645_o;
  /* helpers.vhdl:266:24  */
  assign n3647_o = n3642_o | n3646_o;
  /* helpers.vhdl:266:29  */
  assign n3648_o = n3587_o[21];
  /* helpers.vhdl:266:55  */
  assign n3649_o = n3587_o[20];
  /* helpers.vhdl:266:50  */
  assign n3650_o = ~n3649_o;
  /* helpers.vhdl:266:46  */
  assign n3651_o = n3648_o & n3650_o;
  /* helpers.vhdl:266:24  */
  assign n3652_o = n3647_o | n3651_o;
  /* helpers.vhdl:266:29  */
  assign n3653_o = n3587_o[23];
  /* helpers.vhdl:266:55  */
  assign n3654_o = n3587_o[22];
  /* helpers.vhdl:266:50  */
  assign n3655_o = ~n3654_o;
  /* helpers.vhdl:266:46  */
  assign n3656_o = n3653_o & n3655_o;
  /* helpers.vhdl:266:24  */
  assign n3657_o = n3652_o | n3656_o;
  /* helpers.vhdl:266:29  */
  assign n3658_o = n3587_o[25];
  /* helpers.vhdl:266:55  */
  assign n3659_o = n3587_o[24];
  /* helpers.vhdl:266:50  */
  assign n3660_o = ~n3659_o;
  /* helpers.vhdl:266:46  */
  assign n3661_o = n3658_o & n3660_o;
  /* helpers.vhdl:266:24  */
  assign n3662_o = n3657_o | n3661_o;
  /* helpers.vhdl:266:29  */
  assign n3663_o = n3587_o[27];
  /* helpers.vhdl:266:55  */
  assign n3664_o = n3587_o[26];
  /* helpers.vhdl:266:50  */
  assign n3665_o = ~n3664_o;
  /* helpers.vhdl:266:46  */
  assign n3666_o = n3663_o & n3665_o;
  /* helpers.vhdl:266:24  */
  assign n3667_o = n3662_o | n3666_o;
  /* helpers.vhdl:266:29  */
  assign n3668_o = n3587_o[29];
  /* helpers.vhdl:266:55  */
  assign n3669_o = n3587_o[28];
  /* helpers.vhdl:266:50  */
  assign n3670_o = ~n3669_o;
  /* helpers.vhdl:266:46  */
  assign n3671_o = n3668_o & n3670_o;
  /* helpers.vhdl:266:24  */
  assign n3672_o = n3667_o | n3671_o;
  /* helpers.vhdl:266:29  */
  assign n3673_o = n3587_o[31];
  /* helpers.vhdl:266:55  */
  assign n3674_o = n3587_o[30];
  /* helpers.vhdl:266:50  */
  assign n3675_o = ~n3674_o;
  /* helpers.vhdl:266:46  */
  assign n3676_o = n3673_o & n3675_o;
  /* helpers.vhdl:266:24  */
  assign n3677_o = n3672_o | n3676_o;
  /* helpers.vhdl:266:29  */
  assign n3678_o = n3587_o[33];
  /* helpers.vhdl:266:55  */
  assign n3679_o = n3587_o[32];
  /* helpers.vhdl:266:50  */
  assign n3680_o = ~n3679_o;
  /* helpers.vhdl:266:46  */
  assign n3681_o = n3678_o & n3680_o;
  /* helpers.vhdl:266:24  */
  assign n3682_o = n3677_o | n3681_o;
  /* helpers.vhdl:266:29  */
  assign n3683_o = n3587_o[35];
  /* helpers.vhdl:266:55  */
  assign n3684_o = n3587_o[34];
  /* helpers.vhdl:266:50  */
  assign n3685_o = ~n3684_o;
  /* helpers.vhdl:266:46  */
  assign n3686_o = n3683_o & n3685_o;
  /* helpers.vhdl:266:24  */
  assign n3687_o = n3682_o | n3686_o;
  /* helpers.vhdl:266:29  */
  assign n3688_o = n3587_o[37];
  /* helpers.vhdl:266:55  */
  assign n3689_o = n3587_o[36];
  /* helpers.vhdl:266:50  */
  assign n3690_o = ~n3689_o;
  /* helpers.vhdl:266:46  */
  assign n3691_o = n3688_o & n3690_o;
  /* helpers.vhdl:266:24  */
  assign n3692_o = n3687_o | n3691_o;
  /* helpers.vhdl:266:29  */
  assign n3693_o = n3587_o[39];
  /* helpers.vhdl:266:55  */
  assign n3694_o = n3587_o[38];
  /* helpers.vhdl:266:50  */
  assign n3695_o = ~n3694_o;
  /* helpers.vhdl:266:46  */
  assign n3696_o = n3693_o & n3695_o;
  /* helpers.vhdl:266:24  */
  assign n3697_o = n3692_o | n3696_o;
  /* helpers.vhdl:266:29  */
  assign n3698_o = n3587_o[41];
  /* helpers.vhdl:266:55  */
  assign n3699_o = n3587_o[40];
  /* helpers.vhdl:266:50  */
  assign n3700_o = ~n3699_o;
  /* helpers.vhdl:266:46  */
  assign n3701_o = n3698_o & n3700_o;
  /* helpers.vhdl:266:24  */
  assign n3702_o = n3697_o | n3701_o;
  /* helpers.vhdl:266:29  */
  assign n3703_o = n3587_o[43];
  /* helpers.vhdl:266:55  */
  assign n3704_o = n3587_o[42];
  /* helpers.vhdl:266:50  */
  assign n3705_o = ~n3704_o;
  /* helpers.vhdl:266:46  */
  assign n3706_o = n3703_o & n3705_o;
  /* helpers.vhdl:266:24  */
  assign n3707_o = n3702_o | n3706_o;
  /* helpers.vhdl:266:29  */
  assign n3708_o = n3587_o[45];
  /* helpers.vhdl:266:55  */
  assign n3709_o = n3587_o[44];
  /* helpers.vhdl:266:50  */
  assign n3710_o = ~n3709_o;
  /* helpers.vhdl:266:46  */
  assign n3711_o = n3708_o & n3710_o;
  /* helpers.vhdl:266:24  */
  assign n3712_o = n3707_o | n3711_o;
  /* helpers.vhdl:266:29  */
  assign n3713_o = n3587_o[47];
  /* helpers.vhdl:266:55  */
  assign n3714_o = n3587_o[46];
  /* helpers.vhdl:266:50  */
  assign n3715_o = ~n3714_o;
  /* helpers.vhdl:266:46  */
  assign n3716_o = n3713_o & n3715_o;
  /* helpers.vhdl:266:24  */
  assign n3717_o = n3712_o | n3716_o;
  /* helpers.vhdl:266:29  */
  assign n3718_o = n3587_o[49];
  /* helpers.vhdl:266:55  */
  assign n3719_o = n3587_o[48];
  /* helpers.vhdl:266:50  */
  assign n3720_o = ~n3719_o;
  /* helpers.vhdl:266:46  */
  assign n3721_o = n3718_o & n3720_o;
  /* helpers.vhdl:266:24  */
  assign n3722_o = n3717_o | n3721_o;
  /* helpers.vhdl:266:29  */
  assign n3723_o = n3587_o[51];
  /* helpers.vhdl:266:55  */
  assign n3724_o = n3587_o[50];
  /* helpers.vhdl:266:50  */
  assign n3725_o = ~n3724_o;
  /* helpers.vhdl:266:46  */
  assign n3726_o = n3723_o & n3725_o;
  /* helpers.vhdl:266:24  */
  assign n3727_o = n3722_o | n3726_o;
  /* helpers.vhdl:266:29  */
  assign n3728_o = n3587_o[53];
  /* helpers.vhdl:266:55  */
  assign n3729_o = n3587_o[52];
  /* helpers.vhdl:266:50  */
  assign n3730_o = ~n3729_o;
  /* helpers.vhdl:266:46  */
  assign n3731_o = n3728_o & n3730_o;
  /* helpers.vhdl:266:24  */
  assign n3732_o = n3727_o | n3731_o;
  /* helpers.vhdl:266:29  */
  assign n3733_o = n3587_o[55];
  /* helpers.vhdl:266:55  */
  assign n3734_o = n3587_o[54];
  /* helpers.vhdl:266:50  */
  assign n3735_o = ~n3734_o;
  /* helpers.vhdl:266:46  */
  assign n3736_o = n3733_o & n3735_o;
  /* helpers.vhdl:266:24  */
  assign n3737_o = n3732_o | n3736_o;
  /* helpers.vhdl:266:29  */
  assign n3738_o = n3587_o[57];
  /* helpers.vhdl:266:55  */
  assign n3739_o = n3587_o[56];
  /* helpers.vhdl:266:50  */
  assign n3740_o = ~n3739_o;
  /* helpers.vhdl:266:46  */
  assign n3741_o = n3738_o & n3740_o;
  /* helpers.vhdl:266:24  */
  assign n3742_o = n3737_o | n3741_o;
  /* helpers.vhdl:266:29  */
  assign n3743_o = n3587_o[59];
  /* helpers.vhdl:266:55  */
  assign n3744_o = n3587_o[58];
  /* helpers.vhdl:266:50  */
  assign n3745_o = ~n3744_o;
  /* helpers.vhdl:266:46  */
  assign n3746_o = n3743_o & n3745_o;
  /* helpers.vhdl:266:24  */
  assign n3747_o = n3742_o | n3746_o;
  /* helpers.vhdl:266:29  */
  assign n3748_o = n3587_o[61];
  /* helpers.vhdl:266:55  */
  assign n3749_o = n3587_o[60];
  /* helpers.vhdl:266:50  */
  assign n3750_o = ~n3749_o;
  /* helpers.vhdl:266:46  */
  assign n3751_o = n3748_o & n3750_o;
  /* helpers.vhdl:266:24  */
  assign n3752_o = n3747_o | n3751_o;
  /* helpers.vhdl:266:29  */
  assign n3753_o = n3587_o[63];
  /* helpers.vhdl:266:55  */
  assign n3754_o = n3587_o[62];
  /* helpers.vhdl:266:50  */
  assign n3755_o = ~n3754_o;
  /* helpers.vhdl:266:46  */
  assign n3756_o = n3753_o & n3755_o;
  /* helpers.vhdl:266:24  */
  assign n3757_o = n3752_o | n3756_o;
  /* helpers.vhdl:266:29  */
  assign n3760_o = n3587_o[3];
  /* helpers.vhdl:266:55  */
  assign n3761_o = n3587_o[1];
  /* helpers.vhdl:266:50  */
  assign n3762_o = ~n3761_o;
  /* helpers.vhdl:266:46  */
  assign n3763_o = n3760_o & n3762_o;
  /* helpers.vhdl:266:24  */
  assign n3765_o = 1'b0 | n3763_o;
  /* helpers.vhdl:266:29  */
  assign n3767_o = n3587_o[7];
  /* helpers.vhdl:266:55  */
  assign n3768_o = n3587_o[5];
  /* helpers.vhdl:266:50  */
  assign n3769_o = ~n3768_o;
  /* helpers.vhdl:266:46  */
  assign n3770_o = n3767_o & n3769_o;
  /* helpers.vhdl:266:24  */
  assign n3771_o = n3765_o | n3770_o;
  /* helpers.vhdl:266:29  */
  assign n3772_o = n3587_o[11];
  /* helpers.vhdl:266:55  */
  assign n3773_o = n3587_o[9];
  /* helpers.vhdl:266:50  */
  assign n3774_o = ~n3773_o;
  /* helpers.vhdl:266:46  */
  assign n3775_o = n3772_o & n3774_o;
  /* helpers.vhdl:266:24  */
  assign n3776_o = n3771_o | n3775_o;
  /* helpers.vhdl:266:29  */
  assign n3777_o = n3587_o[15];
  /* helpers.vhdl:266:55  */
  assign n3778_o = n3587_o[13];
  /* helpers.vhdl:266:50  */
  assign n3779_o = ~n3778_o;
  /* helpers.vhdl:266:46  */
  assign n3780_o = n3777_o & n3779_o;
  /* helpers.vhdl:266:24  */
  assign n3781_o = n3776_o | n3780_o;
  /* helpers.vhdl:266:29  */
  assign n3782_o = n3587_o[19];
  /* helpers.vhdl:266:55  */
  assign n3783_o = n3587_o[17];
  /* helpers.vhdl:266:50  */
  assign n3784_o = ~n3783_o;
  /* helpers.vhdl:266:46  */
  assign n3785_o = n3782_o & n3784_o;
  /* helpers.vhdl:266:24  */
  assign n3786_o = n3781_o | n3785_o;
  /* helpers.vhdl:266:29  */
  assign n3787_o = n3587_o[23];
  /* helpers.vhdl:266:55  */
  assign n3788_o = n3587_o[21];
  /* helpers.vhdl:266:50  */
  assign n3789_o = ~n3788_o;
  /* helpers.vhdl:266:46  */
  assign n3790_o = n3787_o & n3789_o;
  /* helpers.vhdl:266:24  */
  assign n3791_o = n3786_o | n3790_o;
  /* helpers.vhdl:266:29  */
  assign n3792_o = n3587_o[27];
  /* helpers.vhdl:266:55  */
  assign n3793_o = n3587_o[25];
  /* helpers.vhdl:266:50  */
  assign n3794_o = ~n3793_o;
  /* helpers.vhdl:266:46  */
  assign n3795_o = n3792_o & n3794_o;
  /* helpers.vhdl:266:24  */
  assign n3796_o = n3791_o | n3795_o;
  /* helpers.vhdl:266:29  */
  assign n3797_o = n3587_o[31];
  /* helpers.vhdl:266:55  */
  assign n3798_o = n3587_o[29];
  /* helpers.vhdl:266:50  */
  assign n3799_o = ~n3798_o;
  /* helpers.vhdl:266:46  */
  assign n3800_o = n3797_o & n3799_o;
  /* helpers.vhdl:266:24  */
  assign n3801_o = n3796_o | n3800_o;
  /* helpers.vhdl:266:29  */
  assign n3802_o = n3587_o[35];
  /* helpers.vhdl:266:55  */
  assign n3803_o = n3587_o[33];
  /* helpers.vhdl:266:50  */
  assign n3804_o = ~n3803_o;
  /* helpers.vhdl:266:46  */
  assign n3805_o = n3802_o & n3804_o;
  /* helpers.vhdl:266:24  */
  assign n3806_o = n3801_o | n3805_o;
  /* helpers.vhdl:266:29  */
  assign n3807_o = n3587_o[39];
  /* helpers.vhdl:266:55  */
  assign n3808_o = n3587_o[37];
  /* helpers.vhdl:266:50  */
  assign n3809_o = ~n3808_o;
  /* helpers.vhdl:266:46  */
  assign n3810_o = n3807_o & n3809_o;
  /* helpers.vhdl:266:24  */
  assign n3811_o = n3806_o | n3810_o;
  /* helpers.vhdl:266:29  */
  assign n3812_o = n3587_o[43];
  /* helpers.vhdl:266:55  */
  assign n3813_o = n3587_o[41];
  /* helpers.vhdl:266:50  */
  assign n3814_o = ~n3813_o;
  /* helpers.vhdl:266:46  */
  assign n3815_o = n3812_o & n3814_o;
  /* helpers.vhdl:266:24  */
  assign n3816_o = n3811_o | n3815_o;
  /* helpers.vhdl:266:29  */
  assign n3817_o = n3587_o[47];
  /* helpers.vhdl:266:55  */
  assign n3818_o = n3587_o[45];
  /* helpers.vhdl:266:50  */
  assign n3819_o = ~n3818_o;
  /* helpers.vhdl:266:46  */
  assign n3820_o = n3817_o & n3819_o;
  /* helpers.vhdl:266:24  */
  assign n3821_o = n3816_o | n3820_o;
  /* helpers.vhdl:266:29  */
  assign n3822_o = n3587_o[51];
  /* helpers.vhdl:266:55  */
  assign n3823_o = n3587_o[49];
  /* helpers.vhdl:266:50  */
  assign n3824_o = ~n3823_o;
  /* helpers.vhdl:266:46  */
  assign n3825_o = n3822_o & n3824_o;
  /* helpers.vhdl:266:24  */
  assign n3826_o = n3821_o | n3825_o;
  /* helpers.vhdl:266:29  */
  assign n3827_o = n3587_o[55];
  /* helpers.vhdl:266:55  */
  assign n3828_o = n3587_o[53];
  /* helpers.vhdl:266:50  */
  assign n3829_o = ~n3828_o;
  /* helpers.vhdl:266:46  */
  assign n3830_o = n3827_o & n3829_o;
  /* helpers.vhdl:266:24  */
  assign n3831_o = n3826_o | n3830_o;
  /* helpers.vhdl:266:29  */
  assign n3832_o = n3587_o[59];
  /* helpers.vhdl:266:55  */
  assign n3833_o = n3587_o[57];
  /* helpers.vhdl:266:50  */
  assign n3834_o = ~n3833_o;
  /* helpers.vhdl:266:46  */
  assign n3835_o = n3832_o & n3834_o;
  /* helpers.vhdl:266:24  */
  assign n3836_o = n3831_o | n3835_o;
  /* helpers.vhdl:266:29  */
  assign n3837_o = n3587_o[63];
  /* helpers.vhdl:266:55  */
  assign n3838_o = n3587_o[61];
  /* helpers.vhdl:266:50  */
  assign n3839_o = ~n3838_o;
  /* helpers.vhdl:266:46  */
  assign n3840_o = n3837_o & n3839_o;
  /* helpers.vhdl:266:24  */
  assign n3841_o = n3836_o | n3840_o;
  /* helpers.vhdl:266:29  */
  assign n3843_o = n3587_o[7];
  /* helpers.vhdl:266:55  */
  assign n3844_o = n3587_o[3];
  /* helpers.vhdl:266:50  */
  assign n3845_o = ~n3844_o;
  /* helpers.vhdl:266:46  */
  assign n3846_o = n3843_o & n3845_o;
  /* helpers.vhdl:266:24  */
  assign n3848_o = 1'b0 | n3846_o;
  /* helpers.vhdl:266:29  */
  assign n3850_o = n3587_o[15];
  /* helpers.vhdl:266:55  */
  assign n3851_o = n3587_o[11];
  /* helpers.vhdl:266:50  */
  assign n3852_o = ~n3851_o;
  /* helpers.vhdl:266:46  */
  assign n3853_o = n3850_o & n3852_o;
  /* helpers.vhdl:266:24  */
  assign n3854_o = n3848_o | n3853_o;
  /* helpers.vhdl:266:29  */
  assign n3855_o = n3587_o[23];
  /* helpers.vhdl:266:55  */
  assign n3856_o = n3587_o[19];
  /* helpers.vhdl:266:50  */
  assign n3857_o = ~n3856_o;
  /* helpers.vhdl:266:46  */
  assign n3858_o = n3855_o & n3857_o;
  /* helpers.vhdl:266:24  */
  assign n3859_o = n3854_o | n3858_o;
  /* helpers.vhdl:266:29  */
  assign n3860_o = n3587_o[31];
  /* helpers.vhdl:266:55  */
  assign n3861_o = n3587_o[27];
  /* helpers.vhdl:266:50  */
  assign n3862_o = ~n3861_o;
  /* helpers.vhdl:266:46  */
  assign n3863_o = n3860_o & n3862_o;
  /* helpers.vhdl:266:24  */
  assign n3864_o = n3859_o | n3863_o;
  /* helpers.vhdl:266:29  */
  assign n3865_o = n3587_o[39];
  /* helpers.vhdl:266:55  */
  assign n3866_o = n3587_o[35];
  /* helpers.vhdl:266:50  */
  assign n3867_o = ~n3866_o;
  /* helpers.vhdl:266:46  */
  assign n3868_o = n3865_o & n3867_o;
  /* helpers.vhdl:266:24  */
  assign n3869_o = n3864_o | n3868_o;
  /* helpers.vhdl:266:29  */
  assign n3870_o = n3587_o[47];
  /* helpers.vhdl:266:55  */
  assign n3871_o = n3587_o[43];
  /* helpers.vhdl:266:50  */
  assign n3872_o = ~n3871_o;
  /* helpers.vhdl:266:46  */
  assign n3873_o = n3870_o & n3872_o;
  /* helpers.vhdl:266:24  */
  assign n3874_o = n3869_o | n3873_o;
  /* helpers.vhdl:266:29  */
  assign n3875_o = n3587_o[55];
  /* helpers.vhdl:266:55  */
  assign n3876_o = n3587_o[51];
  /* helpers.vhdl:266:50  */
  assign n3877_o = ~n3876_o;
  /* helpers.vhdl:266:46  */
  assign n3878_o = n3875_o & n3877_o;
  /* helpers.vhdl:266:24  */
  assign n3879_o = n3874_o | n3878_o;
  /* helpers.vhdl:266:29  */
  assign n3880_o = n3587_o[63];
  /* helpers.vhdl:266:55  */
  assign n3881_o = n3587_o[59];
  /* helpers.vhdl:266:50  */
  assign n3882_o = ~n3881_o;
  /* helpers.vhdl:266:46  */
  assign n3883_o = n3880_o & n3882_o;
  /* helpers.vhdl:266:24  */
  assign n3884_o = n3879_o | n3883_o;
  /* helpers.vhdl:266:29  */
  assign n3886_o = n3587_o[15];
  /* helpers.vhdl:266:55  */
  assign n3887_o = n3587_o[7];
  /* helpers.vhdl:266:50  */
  assign n3888_o = ~n3887_o;
  /* helpers.vhdl:266:46  */
  assign n3889_o = n3886_o & n3888_o;
  /* helpers.vhdl:266:24  */
  assign n3891_o = 1'b0 | n3889_o;
  /* helpers.vhdl:266:29  */
  assign n3893_o = n3587_o[31];
  /* helpers.vhdl:266:55  */
  assign n3894_o = n3587_o[23];
  /* helpers.vhdl:266:50  */
  assign n3895_o = ~n3894_o;
  /* helpers.vhdl:266:46  */
  assign n3896_o = n3893_o & n3895_o;
  /* helpers.vhdl:266:24  */
  assign n3897_o = n3891_o | n3896_o;
  /* helpers.vhdl:266:29  */
  assign n3898_o = n3587_o[47];
  /* helpers.vhdl:266:55  */
  assign n3899_o = n3587_o[39];
  /* helpers.vhdl:266:50  */
  assign n3900_o = ~n3899_o;
  /* helpers.vhdl:266:46  */
  assign n3901_o = n3898_o & n3900_o;
  /* helpers.vhdl:266:24  */
  assign n3902_o = n3897_o | n3901_o;
  /* helpers.vhdl:266:29  */
  assign n3903_o = n3587_o[63];
  /* helpers.vhdl:266:55  */
  assign n3904_o = n3587_o[55];
  /* helpers.vhdl:266:50  */
  assign n3905_o = ~n3904_o;
  /* helpers.vhdl:266:46  */
  assign n3906_o = n3903_o & n3905_o;
  /* helpers.vhdl:266:24  */
  assign n3907_o = n3902_o | n3906_o;
  /* helpers.vhdl:266:29  */
  assign n3909_o = n3587_o[31];
  /* helpers.vhdl:266:55  */
  assign n3910_o = n3587_o[15];
  /* helpers.vhdl:266:50  */
  assign n3911_o = ~n3910_o;
  /* helpers.vhdl:266:46  */
  assign n3912_o = n3909_o & n3911_o;
  /* helpers.vhdl:266:24  */
  assign n3914_o = 1'b0 | n3912_o;
  /* helpers.vhdl:266:29  */
  assign n3916_o = n3587_o[63];
  /* helpers.vhdl:266:55  */
  assign n3917_o = n3587_o[47];
  /* helpers.vhdl:266:50  */
  assign n3918_o = ~n3917_o;
  /* helpers.vhdl:266:46  */
  assign n3919_o = n3916_o & n3918_o;
  /* helpers.vhdl:266:24  */
  assign n3920_o = n3914_o | n3919_o;
  /* helpers.vhdl:266:29  */
  assign n3922_o = n3587_o[63];
  /* helpers.vhdl:266:55  */
  assign n3923_o = n3587_o[31];
  /* helpers.vhdl:266:50  */
  assign n3924_o = ~n3923_o;
  /* helpers.vhdl:266:46  */
  assign n3925_o = n3922_o & n3924_o;
  /* helpers.vhdl:266:24  */
  assign n3927_o = 1'b0 | n3925_o;
  assign n3929_o = {n3927_o, n3920_o, n3907_o, n3884_o, n3841_o, n3757_o};
  /* helpers.vhdl:286:46  */
  assign n3932_o = {56'b0, n3581_o};  //  uext
  /* helpers.vhdl:244:36  */
  assign n3941_o = n3932_o[1];
  /* helpers.vhdl:244:32  */
  assign n3942_o = |(n3941_o);
  /* helpers.vhdl:244:28  */
  assign n3944_o = 1'b0 | n3942_o;
  /* helpers.vhdl:244:36  */
  assign n3946_o = n3932_o[3];
  /* helpers.vhdl:244:32  */
  assign n3947_o = |(n3946_o);
  /* helpers.vhdl:244:28  */
  assign n3948_o = n3944_o | n3947_o;
  /* helpers.vhdl:244:36  */
  assign n3949_o = n3932_o[5];
  /* helpers.vhdl:244:32  */
  assign n3950_o = |(n3949_o);
  /* helpers.vhdl:244:28  */
  assign n3951_o = n3948_o | n3950_o;
  /* helpers.vhdl:244:36  */
  assign n3952_o = n3932_o[7];
  /* helpers.vhdl:244:32  */
  assign n3953_o = |(n3952_o);
  /* helpers.vhdl:244:28  */
  assign n3954_o = n3951_o | n3953_o;
  /* helpers.vhdl:244:36  */
  assign n3955_o = n3932_o[9];
  /* helpers.vhdl:244:32  */
  assign n3956_o = |(n3955_o);
  /* helpers.vhdl:244:28  */
  assign n3957_o = n3954_o | n3956_o;
  /* helpers.vhdl:244:36  */
  assign n3958_o = n3932_o[11];
  /* helpers.vhdl:244:32  */
  assign n3959_o = |(n3958_o);
  /* helpers.vhdl:244:28  */
  assign n3960_o = n3957_o | n3959_o;
  /* helpers.vhdl:244:36  */
  assign n3961_o = n3932_o[13];
  /* helpers.vhdl:244:32  */
  assign n3962_o = |(n3961_o);
  /* helpers.vhdl:244:28  */
  assign n3963_o = n3960_o | n3962_o;
  /* helpers.vhdl:244:36  */
  assign n3964_o = n3932_o[15];
  /* helpers.vhdl:244:32  */
  assign n3965_o = |(n3964_o);
  /* helpers.vhdl:244:28  */
  assign n3966_o = n3963_o | n3965_o;
  /* helpers.vhdl:244:36  */
  assign n3967_o = n3932_o[17];
  /* helpers.vhdl:244:32  */
  assign n3968_o = |(n3967_o);
  /* helpers.vhdl:244:28  */
  assign n3969_o = n3966_o | n3968_o;
  /* helpers.vhdl:244:36  */
  assign n3970_o = n3932_o[19];
  /* helpers.vhdl:244:32  */
  assign n3971_o = |(n3970_o);
  /* helpers.vhdl:244:28  */
  assign n3972_o = n3969_o | n3971_o;
  /* helpers.vhdl:244:36  */
  assign n3973_o = n3932_o[21];
  /* helpers.vhdl:244:32  */
  assign n3974_o = |(n3973_o);
  /* helpers.vhdl:244:28  */
  assign n3975_o = n3972_o | n3974_o;
  /* helpers.vhdl:244:36  */
  assign n3976_o = n3932_o[23];
  /* helpers.vhdl:244:32  */
  assign n3977_o = |(n3976_o);
  /* helpers.vhdl:244:28  */
  assign n3978_o = n3975_o | n3977_o;
  /* helpers.vhdl:244:36  */
  assign n3979_o = n3932_o[25];
  /* helpers.vhdl:244:32  */
  assign n3980_o = |(n3979_o);
  /* helpers.vhdl:244:28  */
  assign n3981_o = n3978_o | n3980_o;
  /* helpers.vhdl:244:36  */
  assign n3982_o = n3932_o[27];
  /* helpers.vhdl:244:32  */
  assign n3983_o = |(n3982_o);
  /* helpers.vhdl:244:28  */
  assign n3984_o = n3981_o | n3983_o;
  /* helpers.vhdl:244:36  */
  assign n3985_o = n3932_o[29];
  /* helpers.vhdl:244:32  */
  assign n3986_o = |(n3985_o);
  /* helpers.vhdl:244:28  */
  assign n3987_o = n3984_o | n3986_o;
  /* helpers.vhdl:244:36  */
  assign n3988_o = n3932_o[31];
  /* helpers.vhdl:244:32  */
  assign n3989_o = |(n3988_o);
  /* helpers.vhdl:244:28  */
  assign n3990_o = n3987_o | n3989_o;
  /* helpers.vhdl:244:36  */
  assign n3991_o = n3932_o[33];
  /* helpers.vhdl:244:32  */
  assign n3992_o = |(n3991_o);
  /* helpers.vhdl:244:28  */
  assign n3993_o = n3990_o | n3992_o;
  /* helpers.vhdl:244:36  */
  assign n3994_o = n3932_o[35];
  /* helpers.vhdl:244:32  */
  assign n3995_o = |(n3994_o);
  /* helpers.vhdl:244:28  */
  assign n3996_o = n3993_o | n3995_o;
  /* helpers.vhdl:244:36  */
  assign n3997_o = n3932_o[37];
  /* helpers.vhdl:244:32  */
  assign n3998_o = |(n3997_o);
  /* helpers.vhdl:244:28  */
  assign n3999_o = n3996_o | n3998_o;
  /* helpers.vhdl:244:36  */
  assign n4000_o = n3932_o[39];
  /* helpers.vhdl:244:32  */
  assign n4001_o = |(n4000_o);
  /* helpers.vhdl:244:28  */
  assign n4002_o = n3999_o | n4001_o;
  /* helpers.vhdl:244:36  */
  assign n4003_o = n3932_o[41];
  /* helpers.vhdl:244:32  */
  assign n4004_o = |(n4003_o);
  /* helpers.vhdl:244:28  */
  assign n4005_o = n4002_o | n4004_o;
  /* helpers.vhdl:244:36  */
  assign n4006_o = n3932_o[43];
  /* helpers.vhdl:244:32  */
  assign n4007_o = |(n4006_o);
  /* helpers.vhdl:244:28  */
  assign n4008_o = n4005_o | n4007_o;
  /* helpers.vhdl:244:36  */
  assign n4009_o = n3932_o[45];
  /* helpers.vhdl:244:32  */
  assign n4010_o = |(n4009_o);
  /* helpers.vhdl:244:28  */
  assign n4011_o = n4008_o | n4010_o;
  /* helpers.vhdl:244:36  */
  assign n4012_o = n3932_o[47];
  /* helpers.vhdl:244:32  */
  assign n4013_o = |(n4012_o);
  /* helpers.vhdl:244:28  */
  assign n4014_o = n4011_o | n4013_o;
  /* helpers.vhdl:244:36  */
  assign n4015_o = n3932_o[49];
  /* helpers.vhdl:244:32  */
  assign n4016_o = |(n4015_o);
  /* helpers.vhdl:244:28  */
  assign n4017_o = n4014_o | n4016_o;
  /* helpers.vhdl:244:36  */
  assign n4018_o = n3932_o[51];
  /* helpers.vhdl:244:32  */
  assign n4019_o = |(n4018_o);
  /* helpers.vhdl:244:28  */
  assign n4020_o = n4017_o | n4019_o;
  /* helpers.vhdl:244:36  */
  assign n4021_o = n3932_o[53];
  /* helpers.vhdl:244:32  */
  assign n4022_o = |(n4021_o);
  /* helpers.vhdl:244:28  */
  assign n4023_o = n4020_o | n4022_o;
  /* helpers.vhdl:244:36  */
  assign n4024_o = n3932_o[55];
  /* helpers.vhdl:244:32  */
  assign n4025_o = |(n4024_o);
  /* helpers.vhdl:244:28  */
  assign n4026_o = n4023_o | n4025_o;
  /* helpers.vhdl:244:36  */
  assign n4027_o = n3932_o[57];
  /* helpers.vhdl:244:32  */
  assign n4028_o = |(n4027_o);
  /* helpers.vhdl:244:28  */
  assign n4029_o = n4026_o | n4028_o;
  /* helpers.vhdl:244:36  */
  assign n4030_o = n3932_o[59];
  /* helpers.vhdl:244:32  */
  assign n4031_o = |(n4030_o);
  /* helpers.vhdl:244:28  */
  assign n4032_o = n4029_o | n4031_o;
  /* helpers.vhdl:244:36  */
  assign n4033_o = n3932_o[61];
  /* helpers.vhdl:244:32  */
  assign n4034_o = |(n4033_o);
  /* helpers.vhdl:244:28  */
  assign n4035_o = n4032_o | n4034_o;
  /* helpers.vhdl:244:36  */
  assign n4036_o = n3932_o[63];
  /* helpers.vhdl:244:32  */
  assign n4037_o = |(n4036_o);
  /* helpers.vhdl:244:28  */
  assign n4038_o = n4035_o | n4037_o;
  /* helpers.vhdl:244:36  */
  assign n4041_o = n3932_o[3:2];
  /* helpers.vhdl:244:32  */
  assign n4042_o = |(n4041_o);
  /* helpers.vhdl:244:28  */
  assign n4044_o = 1'b0 | n4042_o;
  /* helpers.vhdl:244:36  */
  assign n4046_o = n3932_o[7:6];
  /* helpers.vhdl:244:32  */
  assign n4047_o = |(n4046_o);
  /* helpers.vhdl:244:28  */
  assign n4048_o = n4044_o | n4047_o;
  /* helpers.vhdl:244:36  */
  assign n4049_o = n3932_o[11:10];
  /* helpers.vhdl:244:32  */
  assign n4050_o = |(n4049_o);
  /* helpers.vhdl:244:28  */
  assign n4051_o = n4048_o | n4050_o;
  /* helpers.vhdl:244:36  */
  assign n4052_o = n3932_o[15:14];
  /* helpers.vhdl:244:32  */
  assign n4053_o = |(n4052_o);
  /* helpers.vhdl:244:28  */
  assign n4054_o = n4051_o | n4053_o;
  /* helpers.vhdl:244:36  */
  assign n4055_o = n3932_o[19:18];
  /* helpers.vhdl:244:32  */
  assign n4056_o = |(n4055_o);
  /* helpers.vhdl:244:28  */
  assign n4057_o = n4054_o | n4056_o;
  /* helpers.vhdl:244:36  */
  assign n4058_o = n3932_o[23:22];
  /* helpers.vhdl:244:32  */
  assign n4059_o = |(n4058_o);
  /* helpers.vhdl:244:28  */
  assign n4060_o = n4057_o | n4059_o;
  /* helpers.vhdl:244:36  */
  assign n4061_o = n3932_o[27:26];
  /* helpers.vhdl:244:32  */
  assign n4062_o = |(n4061_o);
  /* helpers.vhdl:244:28  */
  assign n4063_o = n4060_o | n4062_o;
  /* helpers.vhdl:244:36  */
  assign n4064_o = n3932_o[31:30];
  /* helpers.vhdl:244:32  */
  assign n4065_o = |(n4064_o);
  /* helpers.vhdl:244:28  */
  assign n4066_o = n4063_o | n4065_o;
  /* helpers.vhdl:244:36  */
  assign n4067_o = n3932_o[35:34];
  /* helpers.vhdl:244:32  */
  assign n4068_o = |(n4067_o);
  /* helpers.vhdl:244:28  */
  assign n4069_o = n4066_o | n4068_o;
  /* helpers.vhdl:244:36  */
  assign n4070_o = n3932_o[39:38];
  /* helpers.vhdl:244:32  */
  assign n4071_o = |(n4070_o);
  /* helpers.vhdl:244:28  */
  assign n4072_o = n4069_o | n4071_o;
  /* helpers.vhdl:244:36  */
  assign n4073_o = n3932_o[43:42];
  /* helpers.vhdl:244:32  */
  assign n4074_o = |(n4073_o);
  /* helpers.vhdl:244:28  */
  assign n4075_o = n4072_o | n4074_o;
  /* helpers.vhdl:244:36  */
  assign n4076_o = n3932_o[47:46];
  /* helpers.vhdl:244:32  */
  assign n4077_o = |(n4076_o);
  /* helpers.vhdl:244:28  */
  assign n4078_o = n4075_o | n4077_o;
  /* helpers.vhdl:244:36  */
  assign n4079_o = n3932_o[51:50];
  /* helpers.vhdl:244:32  */
  assign n4080_o = |(n4079_o);
  /* helpers.vhdl:244:28  */
  assign n4081_o = n4078_o | n4080_o;
  /* helpers.vhdl:244:36  */
  assign n4082_o = n3932_o[55:54];
  /* helpers.vhdl:244:32  */
  assign n4083_o = |(n4082_o);
  /* helpers.vhdl:244:28  */
  assign n4084_o = n4081_o | n4083_o;
  /* helpers.vhdl:244:36  */
  assign n4085_o = n3932_o[59:58];
  /* helpers.vhdl:244:32  */
  assign n4086_o = |(n4085_o);
  /* helpers.vhdl:244:28  */
  assign n4087_o = n4084_o | n4086_o;
  /* helpers.vhdl:244:36  */
  assign n4088_o = n3932_o[63:62];
  /* helpers.vhdl:244:32  */
  assign n4089_o = |(n4088_o);
  /* helpers.vhdl:244:28  */
  assign n4090_o = n4087_o | n4089_o;
  /* helpers.vhdl:244:36  */
  assign n4092_o = n3932_o[7:4];
  /* helpers.vhdl:244:32  */
  assign n4093_o = |(n4092_o);
  /* helpers.vhdl:244:28  */
  assign n4095_o = 1'b0 | n4093_o;
  /* helpers.vhdl:244:36  */
  assign n4097_o = n3932_o[15:12];
  /* helpers.vhdl:244:32  */
  assign n4098_o = |(n4097_o);
  /* helpers.vhdl:244:28  */
  assign n4099_o = n4095_o | n4098_o;
  /* helpers.vhdl:244:36  */
  assign n4100_o = n3932_o[23:20];
  /* helpers.vhdl:244:32  */
  assign n4101_o = |(n4100_o);
  /* helpers.vhdl:244:28  */
  assign n4102_o = n4099_o | n4101_o;
  /* helpers.vhdl:244:36  */
  assign n4103_o = n3932_o[31:28];
  /* helpers.vhdl:244:32  */
  assign n4104_o = |(n4103_o);
  /* helpers.vhdl:244:28  */
  assign n4105_o = n4102_o | n4104_o;
  /* helpers.vhdl:244:36  */
  assign n4106_o = n3932_o[39:36];
  /* helpers.vhdl:244:32  */
  assign n4107_o = |(n4106_o);
  /* helpers.vhdl:244:28  */
  assign n4108_o = n4105_o | n4107_o;
  /* helpers.vhdl:244:36  */
  assign n4109_o = n3932_o[47:44];
  /* helpers.vhdl:244:32  */
  assign n4110_o = |(n4109_o);
  /* helpers.vhdl:244:28  */
  assign n4111_o = n4108_o | n4110_o;
  /* helpers.vhdl:244:36  */
  assign n4112_o = n3932_o[55:52];
  /* helpers.vhdl:244:32  */
  assign n4113_o = |(n4112_o);
  /* helpers.vhdl:244:28  */
  assign n4114_o = n4111_o | n4113_o;
  /* helpers.vhdl:244:36  */
  assign n4115_o = n3932_o[63:60];
  /* helpers.vhdl:244:32  */
  assign n4116_o = |(n4115_o);
  /* helpers.vhdl:244:28  */
  assign n4117_o = n4114_o | n4116_o;
  /* helpers.vhdl:244:36  */
  assign n4119_o = n3932_o[15:8];
  /* helpers.vhdl:244:32  */
  assign n4120_o = |(n4119_o);
  /* helpers.vhdl:244:28  */
  assign n4122_o = 1'b0 | n4120_o;
  /* helpers.vhdl:244:36  */
  assign n4124_o = n3932_o[31:24];
  /* helpers.vhdl:244:32  */
  assign n4125_o = |(n4124_o);
  /* helpers.vhdl:244:28  */
  assign n4126_o = n4122_o | n4125_o;
  /* helpers.vhdl:244:36  */
  assign n4127_o = n3932_o[47:40];
  /* helpers.vhdl:244:32  */
  assign n4128_o = |(n4127_o);
  /* helpers.vhdl:244:28  */
  assign n4129_o = n4126_o | n4128_o;
  /* helpers.vhdl:244:36  */
  assign n4130_o = n3932_o[63:56];
  /* helpers.vhdl:244:32  */
  assign n4131_o = |(n4130_o);
  /* helpers.vhdl:244:28  */
  assign n4132_o = n4129_o | n4131_o;
  /* helpers.vhdl:244:36  */
  assign n4134_o = n3932_o[31:16];
  /* helpers.vhdl:244:32  */
  assign n4135_o = |(n4134_o);
  /* helpers.vhdl:244:28  */
  assign n4137_o = 1'b0 | n4135_o;
  /* helpers.vhdl:244:36  */
  assign n4139_o = n3932_o[63:48];
  /* helpers.vhdl:244:32  */
  assign n4140_o = |(n4139_o);
  /* helpers.vhdl:244:28  */
  assign n4141_o = n4137_o | n4140_o;
  /* helpers.vhdl:244:36  */
  assign n4143_o = n3932_o[63:32];
  /* helpers.vhdl:244:32  */
  assign n4144_o = |(n4143_o);
  /* helpers.vhdl:244:28  */
  assign n4146_o = 1'b0 | n4144_o;
  assign n4148_o = {n4146_o, n4141_o, n4132_o, n4117_o, n4090_o, n4038_o};
  /* helpers.vhdl:287:19  */
  assign n4150_o = n3929_o[5:2];
  /* helpers.vhdl:287:38  */
  assign n4151_o = n4148_o[1:0];
  /* helpers.vhdl:287:32  */
  assign n4152_o = {n4150_o, n4151_o};
  /* xics.vhdl:308:17  */
  assign n4155_o = n4152_o[2:0];
  /* xics.vhdl:440:27  */
  assign n4156_o = int_level_l[0];
  /* xics.vhdl:440:46  */
  assign n4157_o = xives[47:45];
  /* xics.vhdl:440:50  */
  assign n4158_o = n4157_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4159_o = n4158_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4160_o = n4156_o & n4159_o;
  /* xics.vhdl:440:13  */
  assign n4163_o = n4160_o ? 1'b1 : 1'b0;
  /* xics.vhdl:440:27  */
  assign n4166_o = int_level_l[1];
  /* xics.vhdl:440:46  */
  assign n4167_o = xives[44:42];
  /* xics.vhdl:440:50  */
  assign n4168_o = n4167_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4169_o = n4168_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4170_o = n4166_o & n4169_o;
  assign n4172_o = n4164_o[1];
  /* xics.vhdl:440:13  */
  assign n4173_o = n4170_o ? 1'b1 : n4172_o;
  /* xics.vhdl:440:27  */
  assign n4175_o = int_level_l[2];
  /* xics.vhdl:440:46  */
  assign n4176_o = xives[41:39];
  /* xics.vhdl:440:50  */
  assign n4177_o = n4176_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4178_o = n4177_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4179_o = n4175_o & n4178_o;
  assign n4181_o = n4164_o[2];
  /* xics.vhdl:440:13  */
  assign n4182_o = n4179_o ? 1'b1 : n4181_o;
  /* xics.vhdl:440:27  */
  assign n4184_o = int_level_l[3];
  /* xics.vhdl:440:46  */
  assign n4185_o = xives[38:36];
  /* xics.vhdl:440:50  */
  assign n4186_o = n4185_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4187_o = n4186_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4188_o = n4184_o & n4187_o;
  assign n4190_o = n4164_o[3];
  /* xics.vhdl:440:13  */
  assign n4191_o = n4188_o ? 1'b1 : n4190_o;
  /* xics.vhdl:440:27  */
  assign n4193_o = int_level_l[4];
  /* xics.vhdl:440:46  */
  assign n4194_o = xives[35:33];
  /* xics.vhdl:440:50  */
  assign n4195_o = n4194_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4196_o = n4195_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4197_o = n4193_o & n4196_o;
  assign n4199_o = n4164_o[4];
  /* xics.vhdl:440:13  */
  assign n4200_o = n4197_o ? 1'b1 : n4199_o;
  /* xics.vhdl:440:27  */
  assign n4202_o = int_level_l[5];
  /* xics.vhdl:440:46  */
  assign n4203_o = xives[32:30];
  /* xics.vhdl:440:50  */
  assign n4204_o = n4203_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4205_o = n4204_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4206_o = n4202_o & n4205_o;
  assign n4208_o = n4164_o[5];
  /* xics.vhdl:440:13  */
  assign n4209_o = n4206_o ? 1'b1 : n4208_o;
  /* xics.vhdl:440:27  */
  assign n4211_o = int_level_l[6];
  /* xics.vhdl:440:46  */
  assign n4212_o = xives[29:27];
  /* xics.vhdl:440:50  */
  assign n4213_o = n4212_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4214_o = n4213_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4215_o = n4211_o & n4214_o;
  assign n4217_o = n4164_o[6];
  /* xics.vhdl:440:13  */
  assign n4218_o = n4215_o ? 1'b1 : n4217_o;
  /* xics.vhdl:440:27  */
  assign n4220_o = int_level_l[7];
  /* xics.vhdl:440:46  */
  assign n4221_o = xives[26:24];
  /* xics.vhdl:440:50  */
  assign n4222_o = n4221_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4223_o = n4222_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4224_o = n4220_o & n4223_o;
  assign n4226_o = n4164_o[7];
  /* xics.vhdl:440:13  */
  assign n4227_o = n4224_o ? 1'b1 : n4226_o;
  /* xics.vhdl:440:27  */
  assign n4229_o = int_level_l[8];
  /* xics.vhdl:440:46  */
  assign n4230_o = xives[23:21];
  /* xics.vhdl:440:50  */
  assign n4231_o = n4230_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4232_o = n4231_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4233_o = n4229_o & n4232_o;
  assign n4235_o = n4164_o[8];
  /* xics.vhdl:440:13  */
  assign n4236_o = n4233_o ? 1'b1 : n4235_o;
  /* xics.vhdl:440:27  */
  assign n4238_o = int_level_l[9];
  /* xics.vhdl:440:46  */
  assign n4239_o = xives[20:18];
  /* xics.vhdl:440:50  */
  assign n4240_o = n4239_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4241_o = n4240_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4242_o = n4238_o & n4241_o;
  assign n4244_o = n4164_o[9];
  /* xics.vhdl:440:13  */
  assign n4245_o = n4242_o ? 1'b1 : n4244_o;
  /* xics.vhdl:440:27  */
  assign n4247_o = int_level_l[10];
  /* xics.vhdl:440:46  */
  assign n4248_o = xives[17:15];
  /* xics.vhdl:440:50  */
  assign n4249_o = n4248_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4250_o = n4249_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4251_o = n4247_o & n4250_o;
  assign n4253_o = n4164_o[10];
  /* xics.vhdl:440:13  */
  assign n4254_o = n4251_o ? 1'b1 : n4253_o;
  /* xics.vhdl:440:27  */
  assign n4256_o = int_level_l[11];
  /* xics.vhdl:440:46  */
  assign n4257_o = xives[14:12];
  /* xics.vhdl:440:50  */
  assign n4258_o = n4257_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4259_o = n4258_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4260_o = n4256_o & n4259_o;
  assign n4262_o = n4164_o[11];
  /* xics.vhdl:440:13  */
  assign n4263_o = n4260_o ? 1'b1 : n4262_o;
  /* xics.vhdl:440:27  */
  assign n4265_o = int_level_l[12];
  /* xics.vhdl:440:46  */
  assign n4266_o = xives[11:9];
  /* xics.vhdl:440:50  */
  assign n4267_o = n4266_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4268_o = n4267_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4269_o = n4265_o & n4268_o;
  assign n4271_o = n4164_o[12];
  /* xics.vhdl:440:13  */
  assign n4272_o = n4269_o ? 1'b1 : n4271_o;
  /* xics.vhdl:440:27  */
  assign n4274_o = int_level_l[13];
  /* xics.vhdl:440:46  */
  assign n4275_o = xives[8:6];
  /* xics.vhdl:440:50  */
  assign n4276_o = n4275_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4277_o = n4276_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4278_o = n4274_o & n4277_o;
  assign n4280_o = n4164_o[13];
  /* xics.vhdl:440:13  */
  assign n4281_o = n4278_o ? 1'b1 : n4280_o;
  /* xics.vhdl:440:27  */
  assign n4283_o = int_level_l[14];
  /* xics.vhdl:440:46  */
  assign n4284_o = xives[5:3];
  /* xics.vhdl:440:50  */
  assign n4285_o = n4284_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4286_o = n4285_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4287_o = n4283_o & n4286_o;
  assign n4289_o = n4164_o[14];
  /* xics.vhdl:440:13  */
  assign n4290_o = n4287_o ? 1'b1 : n4289_o;
  assign n4291_o = n4164_o[15];
  /* xics.vhdl:440:27  */
  assign n4292_o = int_level_l[15];
  /* xics.vhdl:440:46  */
  assign n4293_o = xives[2:0];
  /* xics.vhdl:440:50  */
  assign n4294_o = n4293_o[2:0];
  /* xics.vhdl:440:54  */
  assign n4295_o = n4294_o == n4155_o;
  /* xics.vhdl:440:37  */
  assign n4296_o = n4292_o & n4295_o;
  /* xics.vhdl:440:13  */
  assign n4298_o = n4296_o ? 1'b1 : n4291_o;
  assign n4306_o = {n4298_o, n4290_o, n4281_o, n4272_o, n4263_o, n4254_o, n4245_o, n4236_o, n4227_o, n4218_o, n4209_o, n4200_o, n4191_o, n4182_o, n4173_o, n4163_o};
  assign n4309_o = n4306_o[14:0];
  assign n4321_o = {1'b1, n4309_o};
  /* helpers.vhdl:282:34  */
  assign n4322_o = -n4321_o;
  assign n4324_o = {1'b1, n4309_o};
  /* helpers.vhdl:283:23  */
  assign n4325_o = n4322_o & n4324_o;
  assign n4327_o = {1'b1, n4309_o};
  /* helpers.vhdl:284:21  */
  assign n4328_o = n4322_o | n4327_o;
  /* helpers.vhdl:285:48  */
  assign n4331_o = {{48{n4328_o[15]}}, n4328_o}; // sext
  /* helpers.vhdl:266:29  */
  assign n4340_o = n4331_o[1];
  /* helpers.vhdl:266:55  */
  assign n4341_o = n4331_o[0];
  /* helpers.vhdl:266:50  */
  assign n4342_o = ~n4341_o;
  /* helpers.vhdl:266:46  */
  assign n4343_o = n4340_o & n4342_o;
  /* helpers.vhdl:266:24  */
  assign n4345_o = 1'b0 | n4343_o;
  /* helpers.vhdl:266:29  */
  assign n4347_o = n4331_o[3];
  /* helpers.vhdl:266:55  */
  assign n4348_o = n4331_o[2];
  /* helpers.vhdl:266:50  */
  assign n4349_o = ~n4348_o;
  /* helpers.vhdl:266:46  */
  assign n4350_o = n4347_o & n4349_o;
  /* helpers.vhdl:266:24  */
  assign n4351_o = n4345_o | n4350_o;
  /* helpers.vhdl:266:29  */
  assign n4352_o = n4331_o[5];
  /* helpers.vhdl:266:55  */
  assign n4353_o = n4331_o[4];
  /* helpers.vhdl:266:50  */
  assign n4354_o = ~n4353_o;
  /* helpers.vhdl:266:46  */
  assign n4355_o = n4352_o & n4354_o;
  /* helpers.vhdl:266:24  */
  assign n4356_o = n4351_o | n4355_o;
  /* helpers.vhdl:266:29  */
  assign n4357_o = n4331_o[7];
  /* helpers.vhdl:266:55  */
  assign n4358_o = n4331_o[6];
  /* helpers.vhdl:266:50  */
  assign n4359_o = ~n4358_o;
  /* helpers.vhdl:266:46  */
  assign n4360_o = n4357_o & n4359_o;
  /* helpers.vhdl:266:24  */
  assign n4361_o = n4356_o | n4360_o;
  /* helpers.vhdl:266:29  */
  assign n4362_o = n4331_o[9];
  /* helpers.vhdl:266:55  */
  assign n4363_o = n4331_o[8];
  /* helpers.vhdl:266:50  */
  assign n4364_o = ~n4363_o;
  /* helpers.vhdl:266:46  */
  assign n4365_o = n4362_o & n4364_o;
  /* helpers.vhdl:266:24  */
  assign n4366_o = n4361_o | n4365_o;
  /* helpers.vhdl:266:29  */
  assign n4367_o = n4331_o[11];
  /* helpers.vhdl:266:55  */
  assign n4368_o = n4331_o[10];
  /* helpers.vhdl:266:50  */
  assign n4369_o = ~n4368_o;
  /* helpers.vhdl:266:46  */
  assign n4370_o = n4367_o & n4369_o;
  /* helpers.vhdl:266:24  */
  assign n4371_o = n4366_o | n4370_o;
  /* helpers.vhdl:266:29  */
  assign n4372_o = n4331_o[13];
  /* helpers.vhdl:266:55  */
  assign n4373_o = n4331_o[12];
  /* helpers.vhdl:266:50  */
  assign n4374_o = ~n4373_o;
  /* helpers.vhdl:266:46  */
  assign n4375_o = n4372_o & n4374_o;
  /* helpers.vhdl:266:24  */
  assign n4376_o = n4371_o | n4375_o;
  /* helpers.vhdl:266:29  */
  assign n4377_o = n4331_o[15];
  /* helpers.vhdl:266:55  */
  assign n4378_o = n4331_o[14];
  /* helpers.vhdl:266:50  */
  assign n4379_o = ~n4378_o;
  /* helpers.vhdl:266:46  */
  assign n4380_o = n4377_o & n4379_o;
  /* helpers.vhdl:266:24  */
  assign n4381_o = n4376_o | n4380_o;
  /* helpers.vhdl:266:29  */
  assign n4382_o = n4331_o[17];
  /* helpers.vhdl:266:55  */
  assign n4383_o = n4331_o[16];
  /* helpers.vhdl:266:50  */
  assign n4384_o = ~n4383_o;
  /* helpers.vhdl:266:46  */
  assign n4385_o = n4382_o & n4384_o;
  /* helpers.vhdl:266:24  */
  assign n4386_o = n4381_o | n4385_o;
  /* helpers.vhdl:266:29  */
  assign n4387_o = n4331_o[19];
  /* helpers.vhdl:266:55  */
  assign n4388_o = n4331_o[18];
  /* helpers.vhdl:266:50  */
  assign n4389_o = ~n4388_o;
  /* helpers.vhdl:266:46  */
  assign n4390_o = n4387_o & n4389_o;
  /* helpers.vhdl:266:24  */
  assign n4391_o = n4386_o | n4390_o;
  /* helpers.vhdl:266:29  */
  assign n4392_o = n4331_o[21];
  /* helpers.vhdl:266:55  */
  assign n4393_o = n4331_o[20];
  /* helpers.vhdl:266:50  */
  assign n4394_o = ~n4393_o;
  /* helpers.vhdl:266:46  */
  assign n4395_o = n4392_o & n4394_o;
  /* helpers.vhdl:266:24  */
  assign n4396_o = n4391_o | n4395_o;
  /* helpers.vhdl:266:29  */
  assign n4397_o = n4331_o[23];
  /* helpers.vhdl:266:55  */
  assign n4398_o = n4331_o[22];
  /* helpers.vhdl:266:50  */
  assign n4399_o = ~n4398_o;
  /* helpers.vhdl:266:46  */
  assign n4400_o = n4397_o & n4399_o;
  /* helpers.vhdl:266:24  */
  assign n4401_o = n4396_o | n4400_o;
  /* helpers.vhdl:266:29  */
  assign n4402_o = n4331_o[25];
  /* helpers.vhdl:266:55  */
  assign n4403_o = n4331_o[24];
  /* helpers.vhdl:266:50  */
  assign n4404_o = ~n4403_o;
  /* helpers.vhdl:266:46  */
  assign n4405_o = n4402_o & n4404_o;
  /* helpers.vhdl:266:24  */
  assign n4406_o = n4401_o | n4405_o;
  /* helpers.vhdl:266:29  */
  assign n4407_o = n4331_o[27];
  /* helpers.vhdl:266:55  */
  assign n4408_o = n4331_o[26];
  /* helpers.vhdl:266:50  */
  assign n4409_o = ~n4408_o;
  /* helpers.vhdl:266:46  */
  assign n4410_o = n4407_o & n4409_o;
  /* helpers.vhdl:266:24  */
  assign n4411_o = n4406_o | n4410_o;
  /* helpers.vhdl:266:29  */
  assign n4412_o = n4331_o[29];
  /* helpers.vhdl:266:55  */
  assign n4413_o = n4331_o[28];
  /* helpers.vhdl:266:50  */
  assign n4414_o = ~n4413_o;
  /* helpers.vhdl:266:46  */
  assign n4415_o = n4412_o & n4414_o;
  /* helpers.vhdl:266:24  */
  assign n4416_o = n4411_o | n4415_o;
  /* helpers.vhdl:266:29  */
  assign n4417_o = n4331_o[31];
  /* helpers.vhdl:266:55  */
  assign n4418_o = n4331_o[30];
  /* helpers.vhdl:266:50  */
  assign n4419_o = ~n4418_o;
  /* helpers.vhdl:266:46  */
  assign n4420_o = n4417_o & n4419_o;
  /* helpers.vhdl:266:24  */
  assign n4421_o = n4416_o | n4420_o;
  /* helpers.vhdl:266:29  */
  assign n4422_o = n4331_o[33];
  /* helpers.vhdl:266:55  */
  assign n4423_o = n4331_o[32];
  /* helpers.vhdl:266:50  */
  assign n4424_o = ~n4423_o;
  /* helpers.vhdl:266:46  */
  assign n4425_o = n4422_o & n4424_o;
  /* helpers.vhdl:266:24  */
  assign n4426_o = n4421_o | n4425_o;
  /* helpers.vhdl:266:29  */
  assign n4427_o = n4331_o[35];
  /* helpers.vhdl:266:55  */
  assign n4428_o = n4331_o[34];
  /* helpers.vhdl:266:50  */
  assign n4429_o = ~n4428_o;
  /* helpers.vhdl:266:46  */
  assign n4430_o = n4427_o & n4429_o;
  /* helpers.vhdl:266:24  */
  assign n4431_o = n4426_o | n4430_o;
  /* helpers.vhdl:266:29  */
  assign n4432_o = n4331_o[37];
  /* helpers.vhdl:266:55  */
  assign n4433_o = n4331_o[36];
  /* helpers.vhdl:266:50  */
  assign n4434_o = ~n4433_o;
  /* helpers.vhdl:266:46  */
  assign n4435_o = n4432_o & n4434_o;
  /* helpers.vhdl:266:24  */
  assign n4436_o = n4431_o | n4435_o;
  /* helpers.vhdl:266:29  */
  assign n4437_o = n4331_o[39];
  /* helpers.vhdl:266:55  */
  assign n4438_o = n4331_o[38];
  /* helpers.vhdl:266:50  */
  assign n4439_o = ~n4438_o;
  /* helpers.vhdl:266:46  */
  assign n4440_o = n4437_o & n4439_o;
  /* helpers.vhdl:266:24  */
  assign n4441_o = n4436_o | n4440_o;
  /* helpers.vhdl:266:29  */
  assign n4442_o = n4331_o[41];
  /* helpers.vhdl:266:55  */
  assign n4443_o = n4331_o[40];
  /* helpers.vhdl:266:50  */
  assign n4444_o = ~n4443_o;
  /* helpers.vhdl:266:46  */
  assign n4445_o = n4442_o & n4444_o;
  /* helpers.vhdl:266:24  */
  assign n4446_o = n4441_o | n4445_o;
  /* helpers.vhdl:266:29  */
  assign n4447_o = n4331_o[43];
  /* helpers.vhdl:266:55  */
  assign n4448_o = n4331_o[42];
  /* helpers.vhdl:266:50  */
  assign n4449_o = ~n4448_o;
  /* helpers.vhdl:266:46  */
  assign n4450_o = n4447_o & n4449_o;
  /* helpers.vhdl:266:24  */
  assign n4451_o = n4446_o | n4450_o;
  /* helpers.vhdl:266:29  */
  assign n4452_o = n4331_o[45];
  /* helpers.vhdl:266:55  */
  assign n4453_o = n4331_o[44];
  /* helpers.vhdl:266:50  */
  assign n4454_o = ~n4453_o;
  /* helpers.vhdl:266:46  */
  assign n4455_o = n4452_o & n4454_o;
  /* helpers.vhdl:266:24  */
  assign n4456_o = n4451_o | n4455_o;
  /* helpers.vhdl:266:29  */
  assign n4457_o = n4331_o[47];
  /* helpers.vhdl:266:55  */
  assign n4458_o = n4331_o[46];
  /* helpers.vhdl:266:50  */
  assign n4459_o = ~n4458_o;
  /* helpers.vhdl:266:46  */
  assign n4460_o = n4457_o & n4459_o;
  /* helpers.vhdl:266:24  */
  assign n4461_o = n4456_o | n4460_o;
  /* helpers.vhdl:266:29  */
  assign n4462_o = n4331_o[49];
  /* helpers.vhdl:266:55  */
  assign n4463_o = n4331_o[48];
  /* helpers.vhdl:266:50  */
  assign n4464_o = ~n4463_o;
  /* helpers.vhdl:266:46  */
  assign n4465_o = n4462_o & n4464_o;
  /* helpers.vhdl:266:24  */
  assign n4466_o = n4461_o | n4465_o;
  /* helpers.vhdl:266:29  */
  assign n4467_o = n4331_o[51];
  /* helpers.vhdl:266:55  */
  assign n4468_o = n4331_o[50];
  /* helpers.vhdl:266:50  */
  assign n4469_o = ~n4468_o;
  /* helpers.vhdl:266:46  */
  assign n4470_o = n4467_o & n4469_o;
  /* helpers.vhdl:266:24  */
  assign n4471_o = n4466_o | n4470_o;
  /* helpers.vhdl:266:29  */
  assign n4472_o = n4331_o[53];
  /* helpers.vhdl:266:55  */
  assign n4473_o = n4331_o[52];
  /* helpers.vhdl:266:50  */
  assign n4474_o = ~n4473_o;
  /* helpers.vhdl:266:46  */
  assign n4475_o = n4472_o & n4474_o;
  /* helpers.vhdl:266:24  */
  assign n4476_o = n4471_o | n4475_o;
  /* helpers.vhdl:266:29  */
  assign n4477_o = n4331_o[55];
  /* helpers.vhdl:266:55  */
  assign n4478_o = n4331_o[54];
  /* helpers.vhdl:266:50  */
  assign n4479_o = ~n4478_o;
  /* helpers.vhdl:266:46  */
  assign n4480_o = n4477_o & n4479_o;
  /* helpers.vhdl:266:24  */
  assign n4481_o = n4476_o | n4480_o;
  /* helpers.vhdl:266:29  */
  assign n4482_o = n4331_o[57];
  /* helpers.vhdl:266:55  */
  assign n4483_o = n4331_o[56];
  /* helpers.vhdl:266:50  */
  assign n4484_o = ~n4483_o;
  /* helpers.vhdl:266:46  */
  assign n4485_o = n4482_o & n4484_o;
  /* helpers.vhdl:266:24  */
  assign n4486_o = n4481_o | n4485_o;
  /* helpers.vhdl:266:29  */
  assign n4487_o = n4331_o[59];
  /* helpers.vhdl:266:55  */
  assign n4488_o = n4331_o[58];
  /* helpers.vhdl:266:50  */
  assign n4489_o = ~n4488_o;
  /* helpers.vhdl:266:46  */
  assign n4490_o = n4487_o & n4489_o;
  /* helpers.vhdl:266:24  */
  assign n4491_o = n4486_o | n4490_o;
  /* helpers.vhdl:266:29  */
  assign n4492_o = n4331_o[61];
  /* helpers.vhdl:266:55  */
  assign n4493_o = n4331_o[60];
  /* helpers.vhdl:266:50  */
  assign n4494_o = ~n4493_o;
  /* helpers.vhdl:266:46  */
  assign n4495_o = n4492_o & n4494_o;
  /* helpers.vhdl:266:24  */
  assign n4496_o = n4491_o | n4495_o;
  /* helpers.vhdl:266:29  */
  assign n4497_o = n4331_o[63];
  /* helpers.vhdl:266:55  */
  assign n4498_o = n4331_o[62];
  /* helpers.vhdl:266:50  */
  assign n4499_o = ~n4498_o;
  /* helpers.vhdl:266:46  */
  assign n4500_o = n4497_o & n4499_o;
  /* helpers.vhdl:266:24  */
  assign n4501_o = n4496_o | n4500_o;
  /* helpers.vhdl:266:29  */
  assign n4504_o = n4331_o[3];
  /* helpers.vhdl:266:55  */
  assign n4505_o = n4331_o[1];
  /* helpers.vhdl:266:50  */
  assign n4506_o = ~n4505_o;
  /* helpers.vhdl:266:46  */
  assign n4507_o = n4504_o & n4506_o;
  /* helpers.vhdl:266:24  */
  assign n4509_o = 1'b0 | n4507_o;
  /* helpers.vhdl:266:29  */
  assign n4511_o = n4331_o[7];
  /* helpers.vhdl:266:55  */
  assign n4512_o = n4331_o[5];
  /* helpers.vhdl:266:50  */
  assign n4513_o = ~n4512_o;
  /* helpers.vhdl:266:46  */
  assign n4514_o = n4511_o & n4513_o;
  /* helpers.vhdl:266:24  */
  assign n4515_o = n4509_o | n4514_o;
  /* helpers.vhdl:266:29  */
  assign n4516_o = n4331_o[11];
  /* helpers.vhdl:266:55  */
  assign n4517_o = n4331_o[9];
  /* helpers.vhdl:266:50  */
  assign n4518_o = ~n4517_o;
  /* helpers.vhdl:266:46  */
  assign n4519_o = n4516_o & n4518_o;
  /* helpers.vhdl:266:24  */
  assign n4520_o = n4515_o | n4519_o;
  /* helpers.vhdl:266:29  */
  assign n4521_o = n4331_o[15];
  /* helpers.vhdl:266:55  */
  assign n4522_o = n4331_o[13];
  /* helpers.vhdl:266:50  */
  assign n4523_o = ~n4522_o;
  /* helpers.vhdl:266:46  */
  assign n4524_o = n4521_o & n4523_o;
  /* helpers.vhdl:266:24  */
  assign n4525_o = n4520_o | n4524_o;
  /* helpers.vhdl:266:29  */
  assign n4526_o = n4331_o[19];
  /* helpers.vhdl:266:55  */
  assign n4527_o = n4331_o[17];
  /* helpers.vhdl:266:50  */
  assign n4528_o = ~n4527_o;
  /* helpers.vhdl:266:46  */
  assign n4529_o = n4526_o & n4528_o;
  /* helpers.vhdl:266:24  */
  assign n4530_o = n4525_o | n4529_o;
  /* helpers.vhdl:266:29  */
  assign n4531_o = n4331_o[23];
  /* helpers.vhdl:266:55  */
  assign n4532_o = n4331_o[21];
  /* helpers.vhdl:266:50  */
  assign n4533_o = ~n4532_o;
  /* helpers.vhdl:266:46  */
  assign n4534_o = n4531_o & n4533_o;
  /* helpers.vhdl:266:24  */
  assign n4535_o = n4530_o | n4534_o;
  /* helpers.vhdl:266:29  */
  assign n4536_o = n4331_o[27];
  /* helpers.vhdl:266:55  */
  assign n4537_o = n4331_o[25];
  /* helpers.vhdl:266:50  */
  assign n4538_o = ~n4537_o;
  /* helpers.vhdl:266:46  */
  assign n4539_o = n4536_o & n4538_o;
  /* helpers.vhdl:266:24  */
  assign n4540_o = n4535_o | n4539_o;
  /* helpers.vhdl:266:29  */
  assign n4541_o = n4331_o[31];
  /* helpers.vhdl:266:55  */
  assign n4542_o = n4331_o[29];
  /* helpers.vhdl:266:50  */
  assign n4543_o = ~n4542_o;
  /* helpers.vhdl:266:46  */
  assign n4544_o = n4541_o & n4543_o;
  /* helpers.vhdl:266:24  */
  assign n4545_o = n4540_o | n4544_o;
  /* helpers.vhdl:266:29  */
  assign n4546_o = n4331_o[35];
  /* helpers.vhdl:266:55  */
  assign n4547_o = n4331_o[33];
  /* helpers.vhdl:266:50  */
  assign n4548_o = ~n4547_o;
  /* helpers.vhdl:266:46  */
  assign n4549_o = n4546_o & n4548_o;
  /* helpers.vhdl:266:24  */
  assign n4550_o = n4545_o | n4549_o;
  /* helpers.vhdl:266:29  */
  assign n4551_o = n4331_o[39];
  /* helpers.vhdl:266:55  */
  assign n4552_o = n4331_o[37];
  /* helpers.vhdl:266:50  */
  assign n4553_o = ~n4552_o;
  /* helpers.vhdl:266:46  */
  assign n4554_o = n4551_o & n4553_o;
  /* helpers.vhdl:266:24  */
  assign n4555_o = n4550_o | n4554_o;
  /* helpers.vhdl:266:29  */
  assign n4556_o = n4331_o[43];
  /* helpers.vhdl:266:55  */
  assign n4557_o = n4331_o[41];
  /* helpers.vhdl:266:50  */
  assign n4558_o = ~n4557_o;
  /* helpers.vhdl:266:46  */
  assign n4559_o = n4556_o & n4558_o;
  /* helpers.vhdl:266:24  */
  assign n4560_o = n4555_o | n4559_o;
  /* helpers.vhdl:266:29  */
  assign n4561_o = n4331_o[47];
  /* helpers.vhdl:266:55  */
  assign n4562_o = n4331_o[45];
  /* helpers.vhdl:266:50  */
  assign n4563_o = ~n4562_o;
  /* helpers.vhdl:266:46  */
  assign n4564_o = n4561_o & n4563_o;
  /* helpers.vhdl:266:24  */
  assign n4565_o = n4560_o | n4564_o;
  /* helpers.vhdl:266:29  */
  assign n4566_o = n4331_o[51];
  /* helpers.vhdl:266:55  */
  assign n4567_o = n4331_o[49];
  /* helpers.vhdl:266:50  */
  assign n4568_o = ~n4567_o;
  /* helpers.vhdl:266:46  */
  assign n4569_o = n4566_o & n4568_o;
  /* helpers.vhdl:266:24  */
  assign n4570_o = n4565_o | n4569_o;
  /* helpers.vhdl:266:29  */
  assign n4571_o = n4331_o[55];
  /* helpers.vhdl:266:55  */
  assign n4572_o = n4331_o[53];
  /* helpers.vhdl:266:50  */
  assign n4573_o = ~n4572_o;
  /* helpers.vhdl:266:46  */
  assign n4574_o = n4571_o & n4573_o;
  /* helpers.vhdl:266:24  */
  assign n4575_o = n4570_o | n4574_o;
  /* helpers.vhdl:266:29  */
  assign n4576_o = n4331_o[59];
  /* helpers.vhdl:266:55  */
  assign n4577_o = n4331_o[57];
  /* helpers.vhdl:266:50  */
  assign n4578_o = ~n4577_o;
  /* helpers.vhdl:266:46  */
  assign n4579_o = n4576_o & n4578_o;
  /* helpers.vhdl:266:24  */
  assign n4580_o = n4575_o | n4579_o;
  /* helpers.vhdl:266:29  */
  assign n4581_o = n4331_o[63];
  /* helpers.vhdl:266:55  */
  assign n4582_o = n4331_o[61];
  /* helpers.vhdl:266:50  */
  assign n4583_o = ~n4582_o;
  /* helpers.vhdl:266:46  */
  assign n4584_o = n4581_o & n4583_o;
  /* helpers.vhdl:266:24  */
  assign n4585_o = n4580_o | n4584_o;
  /* helpers.vhdl:266:29  */
  assign n4587_o = n4331_o[7];
  /* helpers.vhdl:266:55  */
  assign n4588_o = n4331_o[3];
  /* helpers.vhdl:266:50  */
  assign n4589_o = ~n4588_o;
  /* helpers.vhdl:266:46  */
  assign n4590_o = n4587_o & n4589_o;
  /* helpers.vhdl:266:24  */
  assign n4592_o = 1'b0 | n4590_o;
  /* helpers.vhdl:266:29  */
  assign n4594_o = n4331_o[15];
  /* helpers.vhdl:266:55  */
  assign n4595_o = n4331_o[11];
  /* helpers.vhdl:266:50  */
  assign n4596_o = ~n4595_o;
  /* helpers.vhdl:266:46  */
  assign n4597_o = n4594_o & n4596_o;
  /* helpers.vhdl:266:24  */
  assign n4598_o = n4592_o | n4597_o;
  /* helpers.vhdl:266:29  */
  assign n4599_o = n4331_o[23];
  /* helpers.vhdl:266:55  */
  assign n4600_o = n4331_o[19];
  /* helpers.vhdl:266:50  */
  assign n4601_o = ~n4600_o;
  /* helpers.vhdl:266:46  */
  assign n4602_o = n4599_o & n4601_o;
  /* helpers.vhdl:266:24  */
  assign n4603_o = n4598_o | n4602_o;
  /* helpers.vhdl:266:29  */
  assign n4604_o = n4331_o[31];
  /* helpers.vhdl:266:55  */
  assign n4605_o = n4331_o[27];
  /* helpers.vhdl:266:50  */
  assign n4606_o = ~n4605_o;
  /* helpers.vhdl:266:46  */
  assign n4607_o = n4604_o & n4606_o;
  /* helpers.vhdl:266:24  */
  assign n4608_o = n4603_o | n4607_o;
  /* helpers.vhdl:266:29  */
  assign n4609_o = n4331_o[39];
  /* helpers.vhdl:266:55  */
  assign n4610_o = n4331_o[35];
  /* helpers.vhdl:266:50  */
  assign n4611_o = ~n4610_o;
  /* helpers.vhdl:266:46  */
  assign n4612_o = n4609_o & n4611_o;
  /* helpers.vhdl:266:24  */
  assign n4613_o = n4608_o | n4612_o;
  /* helpers.vhdl:266:29  */
  assign n4614_o = n4331_o[47];
  /* helpers.vhdl:266:55  */
  assign n4615_o = n4331_o[43];
  /* helpers.vhdl:266:50  */
  assign n4616_o = ~n4615_o;
  /* helpers.vhdl:266:46  */
  assign n4617_o = n4614_o & n4616_o;
  /* helpers.vhdl:266:24  */
  assign n4618_o = n4613_o | n4617_o;
  /* helpers.vhdl:266:29  */
  assign n4619_o = n4331_o[55];
  /* helpers.vhdl:266:55  */
  assign n4620_o = n4331_o[51];
  /* helpers.vhdl:266:50  */
  assign n4621_o = ~n4620_o;
  /* helpers.vhdl:266:46  */
  assign n4622_o = n4619_o & n4621_o;
  /* helpers.vhdl:266:24  */
  assign n4623_o = n4618_o | n4622_o;
  /* helpers.vhdl:266:29  */
  assign n4624_o = n4331_o[63];
  /* helpers.vhdl:266:55  */
  assign n4625_o = n4331_o[59];
  /* helpers.vhdl:266:50  */
  assign n4626_o = ~n4625_o;
  /* helpers.vhdl:266:46  */
  assign n4627_o = n4624_o & n4626_o;
  /* helpers.vhdl:266:24  */
  assign n4628_o = n4623_o | n4627_o;
  /* helpers.vhdl:266:29  */
  assign n4630_o = n4331_o[15];
  /* helpers.vhdl:266:55  */
  assign n4631_o = n4331_o[7];
  /* helpers.vhdl:266:50  */
  assign n4632_o = ~n4631_o;
  /* helpers.vhdl:266:46  */
  assign n4633_o = n4630_o & n4632_o;
  /* helpers.vhdl:266:24  */
  assign n4635_o = 1'b0 | n4633_o;
  /* helpers.vhdl:266:29  */
  assign n4637_o = n4331_o[31];
  /* helpers.vhdl:266:55  */
  assign n4638_o = n4331_o[23];
  /* helpers.vhdl:266:50  */
  assign n4639_o = ~n4638_o;
  /* helpers.vhdl:266:46  */
  assign n4640_o = n4637_o & n4639_o;
  /* helpers.vhdl:266:24  */
  assign n4641_o = n4635_o | n4640_o;
  /* helpers.vhdl:266:29  */
  assign n4642_o = n4331_o[47];
  /* helpers.vhdl:266:55  */
  assign n4643_o = n4331_o[39];
  /* helpers.vhdl:266:50  */
  assign n4644_o = ~n4643_o;
  /* helpers.vhdl:266:46  */
  assign n4645_o = n4642_o & n4644_o;
  /* helpers.vhdl:266:24  */
  assign n4646_o = n4641_o | n4645_o;
  /* helpers.vhdl:266:29  */
  assign n4647_o = n4331_o[63];
  /* helpers.vhdl:266:55  */
  assign n4648_o = n4331_o[55];
  /* helpers.vhdl:266:50  */
  assign n4649_o = ~n4648_o;
  /* helpers.vhdl:266:46  */
  assign n4650_o = n4647_o & n4649_o;
  /* helpers.vhdl:266:24  */
  assign n4651_o = n4646_o | n4650_o;
  /* helpers.vhdl:266:29  */
  assign n4653_o = n4331_o[31];
  /* helpers.vhdl:266:55  */
  assign n4654_o = n4331_o[15];
  /* helpers.vhdl:266:50  */
  assign n4655_o = ~n4654_o;
  /* helpers.vhdl:266:46  */
  assign n4656_o = n4653_o & n4655_o;
  /* helpers.vhdl:266:24  */
  assign n4658_o = 1'b0 | n4656_o;
  /* helpers.vhdl:266:29  */
  assign n4660_o = n4331_o[63];
  /* helpers.vhdl:266:55  */
  assign n4661_o = n4331_o[47];
  /* helpers.vhdl:266:50  */
  assign n4662_o = ~n4661_o;
  /* helpers.vhdl:266:46  */
  assign n4663_o = n4660_o & n4662_o;
  /* helpers.vhdl:266:24  */
  assign n4664_o = n4658_o | n4663_o;
  /* helpers.vhdl:266:29  */
  assign n4666_o = n4331_o[63];
  /* helpers.vhdl:266:55  */
  assign n4667_o = n4331_o[31];
  /* helpers.vhdl:266:50  */
  assign n4668_o = ~n4667_o;
  /* helpers.vhdl:266:46  */
  assign n4669_o = n4666_o & n4668_o;
  /* helpers.vhdl:266:24  */
  assign n4671_o = 1'b0 | n4669_o;
  assign n4673_o = {n4671_o, n4664_o, n4651_o, n4628_o, n4585_o, n4501_o};
  /* helpers.vhdl:286:46  */
  assign n4676_o = {48'b0, n4325_o};  //  uext
  /* helpers.vhdl:244:36  */
  assign n4685_o = n4676_o[1];
  /* helpers.vhdl:244:32  */
  assign n4686_o = |(n4685_o);
  /* helpers.vhdl:244:28  */
  assign n4688_o = 1'b0 | n4686_o;
  /* helpers.vhdl:244:36  */
  assign n4690_o = n4676_o[3];
  /* helpers.vhdl:244:32  */
  assign n4691_o = |(n4690_o);
  /* helpers.vhdl:244:28  */
  assign n4692_o = n4688_o | n4691_o;
  /* helpers.vhdl:244:36  */
  assign n4693_o = n4676_o[5];
  /* helpers.vhdl:244:32  */
  assign n4694_o = |(n4693_o);
  /* helpers.vhdl:244:28  */
  assign n4695_o = n4692_o | n4694_o;
  /* helpers.vhdl:244:36  */
  assign n4696_o = n4676_o[7];
  /* helpers.vhdl:244:32  */
  assign n4697_o = |(n4696_o);
  /* helpers.vhdl:244:28  */
  assign n4698_o = n4695_o | n4697_o;
  /* helpers.vhdl:244:36  */
  assign n4699_o = n4676_o[9];
  /* helpers.vhdl:244:32  */
  assign n4700_o = |(n4699_o);
  /* helpers.vhdl:244:28  */
  assign n4701_o = n4698_o | n4700_o;
  /* helpers.vhdl:244:36  */
  assign n4702_o = n4676_o[11];
  /* helpers.vhdl:244:32  */
  assign n4703_o = |(n4702_o);
  /* helpers.vhdl:244:28  */
  assign n4704_o = n4701_o | n4703_o;
  /* helpers.vhdl:244:36  */
  assign n4705_o = n4676_o[13];
  /* helpers.vhdl:244:32  */
  assign n4706_o = |(n4705_o);
  /* helpers.vhdl:244:28  */
  assign n4707_o = n4704_o | n4706_o;
  /* helpers.vhdl:244:36  */
  assign n4708_o = n4676_o[15];
  /* helpers.vhdl:244:32  */
  assign n4709_o = |(n4708_o);
  /* helpers.vhdl:244:28  */
  assign n4710_o = n4707_o | n4709_o;
  /* helpers.vhdl:244:36  */
  assign n4711_o = n4676_o[17];
  /* helpers.vhdl:244:32  */
  assign n4712_o = |(n4711_o);
  /* helpers.vhdl:244:28  */
  assign n4713_o = n4710_o | n4712_o;
  /* helpers.vhdl:244:36  */
  assign n4714_o = n4676_o[19];
  /* helpers.vhdl:244:32  */
  assign n4715_o = |(n4714_o);
  /* helpers.vhdl:244:28  */
  assign n4716_o = n4713_o | n4715_o;
  /* helpers.vhdl:244:36  */
  assign n4717_o = n4676_o[21];
  /* helpers.vhdl:244:32  */
  assign n4718_o = |(n4717_o);
  /* helpers.vhdl:244:28  */
  assign n4719_o = n4716_o | n4718_o;
  /* helpers.vhdl:244:36  */
  assign n4720_o = n4676_o[23];
  /* helpers.vhdl:244:32  */
  assign n4721_o = |(n4720_o);
  /* helpers.vhdl:244:28  */
  assign n4722_o = n4719_o | n4721_o;
  /* helpers.vhdl:244:36  */
  assign n4723_o = n4676_o[25];
  /* helpers.vhdl:244:32  */
  assign n4724_o = |(n4723_o);
  /* helpers.vhdl:244:28  */
  assign n4725_o = n4722_o | n4724_o;
  /* helpers.vhdl:244:36  */
  assign n4726_o = n4676_o[27];
  /* helpers.vhdl:244:32  */
  assign n4727_o = |(n4726_o);
  /* helpers.vhdl:244:28  */
  assign n4728_o = n4725_o | n4727_o;
  /* helpers.vhdl:244:36  */
  assign n4729_o = n4676_o[29];
  /* helpers.vhdl:244:32  */
  assign n4730_o = |(n4729_o);
  /* helpers.vhdl:244:28  */
  assign n4731_o = n4728_o | n4730_o;
  /* helpers.vhdl:244:36  */
  assign n4732_o = n4676_o[31];
  /* helpers.vhdl:244:32  */
  assign n4733_o = |(n4732_o);
  /* helpers.vhdl:244:28  */
  assign n4734_o = n4731_o | n4733_o;
  /* helpers.vhdl:244:36  */
  assign n4735_o = n4676_o[33];
  /* helpers.vhdl:244:32  */
  assign n4736_o = |(n4735_o);
  /* helpers.vhdl:244:28  */
  assign n4737_o = n4734_o | n4736_o;
  /* helpers.vhdl:244:36  */
  assign n4738_o = n4676_o[35];
  /* helpers.vhdl:244:32  */
  assign n4739_o = |(n4738_o);
  /* helpers.vhdl:244:28  */
  assign n4740_o = n4737_o | n4739_o;
  /* helpers.vhdl:244:36  */
  assign n4741_o = n4676_o[37];
  /* helpers.vhdl:244:32  */
  assign n4742_o = |(n4741_o);
  /* helpers.vhdl:244:28  */
  assign n4743_o = n4740_o | n4742_o;
  /* helpers.vhdl:244:36  */
  assign n4744_o = n4676_o[39];
  /* helpers.vhdl:244:32  */
  assign n4745_o = |(n4744_o);
  /* helpers.vhdl:244:28  */
  assign n4746_o = n4743_o | n4745_o;
  /* helpers.vhdl:244:36  */
  assign n4747_o = n4676_o[41];
  /* helpers.vhdl:244:32  */
  assign n4748_o = |(n4747_o);
  /* helpers.vhdl:244:28  */
  assign n4749_o = n4746_o | n4748_o;
  /* helpers.vhdl:244:36  */
  assign n4750_o = n4676_o[43];
  /* helpers.vhdl:244:32  */
  assign n4751_o = |(n4750_o);
  /* helpers.vhdl:244:28  */
  assign n4752_o = n4749_o | n4751_o;
  /* helpers.vhdl:244:36  */
  assign n4753_o = n4676_o[45];
  /* helpers.vhdl:244:32  */
  assign n4754_o = |(n4753_o);
  /* helpers.vhdl:244:28  */
  assign n4755_o = n4752_o | n4754_o;
  /* helpers.vhdl:244:36  */
  assign n4756_o = n4676_o[47];
  /* helpers.vhdl:244:32  */
  assign n4757_o = |(n4756_o);
  /* helpers.vhdl:244:28  */
  assign n4758_o = n4755_o | n4757_o;
  /* helpers.vhdl:244:36  */
  assign n4759_o = n4676_o[49];
  /* helpers.vhdl:244:32  */
  assign n4760_o = |(n4759_o);
  /* helpers.vhdl:244:28  */
  assign n4761_o = n4758_o | n4760_o;
  /* helpers.vhdl:244:36  */
  assign n4762_o = n4676_o[51];
  /* helpers.vhdl:244:32  */
  assign n4763_o = |(n4762_o);
  /* helpers.vhdl:244:28  */
  assign n4764_o = n4761_o | n4763_o;
  /* helpers.vhdl:244:36  */
  assign n4765_o = n4676_o[53];
  /* helpers.vhdl:244:32  */
  assign n4766_o = |(n4765_o);
  /* helpers.vhdl:244:28  */
  assign n4767_o = n4764_o | n4766_o;
  /* helpers.vhdl:244:36  */
  assign n4768_o = n4676_o[55];
  /* helpers.vhdl:244:32  */
  assign n4769_o = |(n4768_o);
  /* helpers.vhdl:244:28  */
  assign n4770_o = n4767_o | n4769_o;
  /* helpers.vhdl:244:36  */
  assign n4771_o = n4676_o[57];
  /* helpers.vhdl:244:32  */
  assign n4772_o = |(n4771_o);
  /* helpers.vhdl:244:28  */
  assign n4773_o = n4770_o | n4772_o;
  /* helpers.vhdl:244:36  */
  assign n4774_o = n4676_o[59];
  /* helpers.vhdl:244:32  */
  assign n4775_o = |(n4774_o);
  /* helpers.vhdl:244:28  */
  assign n4776_o = n4773_o | n4775_o;
  /* helpers.vhdl:244:36  */
  assign n4777_o = n4676_o[61];
  /* helpers.vhdl:244:32  */
  assign n4778_o = |(n4777_o);
  /* helpers.vhdl:244:28  */
  assign n4779_o = n4776_o | n4778_o;
  /* helpers.vhdl:244:36  */
  assign n4780_o = n4676_o[63];
  /* helpers.vhdl:244:32  */
  assign n4781_o = |(n4780_o);
  /* helpers.vhdl:244:28  */
  assign n4782_o = n4779_o | n4781_o;
  /* helpers.vhdl:244:36  */
  assign n4785_o = n4676_o[3:2];
  /* helpers.vhdl:244:32  */
  assign n4786_o = |(n4785_o);
  /* helpers.vhdl:244:28  */
  assign n4788_o = 1'b0 | n4786_o;
  /* helpers.vhdl:244:36  */
  assign n4790_o = n4676_o[7:6];
  /* helpers.vhdl:244:32  */
  assign n4791_o = |(n4790_o);
  /* helpers.vhdl:244:28  */
  assign n4792_o = n4788_o | n4791_o;
  /* helpers.vhdl:244:36  */
  assign n4793_o = n4676_o[11:10];
  /* helpers.vhdl:244:32  */
  assign n4794_o = |(n4793_o);
  /* helpers.vhdl:244:28  */
  assign n4795_o = n4792_o | n4794_o;
  /* helpers.vhdl:244:36  */
  assign n4796_o = n4676_o[15:14];
  /* helpers.vhdl:244:32  */
  assign n4797_o = |(n4796_o);
  /* helpers.vhdl:244:28  */
  assign n4798_o = n4795_o | n4797_o;
  /* helpers.vhdl:244:36  */
  assign n4799_o = n4676_o[19:18];
  /* helpers.vhdl:244:32  */
  assign n4800_o = |(n4799_o);
  /* helpers.vhdl:244:28  */
  assign n4801_o = n4798_o | n4800_o;
  /* helpers.vhdl:244:36  */
  assign n4802_o = n4676_o[23:22];
  /* helpers.vhdl:244:32  */
  assign n4803_o = |(n4802_o);
  /* helpers.vhdl:244:28  */
  assign n4804_o = n4801_o | n4803_o;
  /* helpers.vhdl:244:36  */
  assign n4805_o = n4676_o[27:26];
  /* helpers.vhdl:244:32  */
  assign n4806_o = |(n4805_o);
  /* helpers.vhdl:244:28  */
  assign n4807_o = n4804_o | n4806_o;
  /* helpers.vhdl:244:36  */
  assign n4808_o = n4676_o[31:30];
  /* helpers.vhdl:244:32  */
  assign n4809_o = |(n4808_o);
  /* helpers.vhdl:244:28  */
  assign n4810_o = n4807_o | n4809_o;
  /* helpers.vhdl:244:36  */
  assign n4811_o = n4676_o[35:34];
  /* helpers.vhdl:244:32  */
  assign n4812_o = |(n4811_o);
  /* helpers.vhdl:244:28  */
  assign n4813_o = n4810_o | n4812_o;
  /* helpers.vhdl:244:36  */
  assign n4814_o = n4676_o[39:38];
  /* helpers.vhdl:244:32  */
  assign n4815_o = |(n4814_o);
  /* helpers.vhdl:244:28  */
  assign n4816_o = n4813_o | n4815_o;
  /* helpers.vhdl:244:36  */
  assign n4817_o = n4676_o[43:42];
  /* helpers.vhdl:244:32  */
  assign n4818_o = |(n4817_o);
  /* helpers.vhdl:244:28  */
  assign n4819_o = n4816_o | n4818_o;
  /* helpers.vhdl:244:36  */
  assign n4820_o = n4676_o[47:46];
  /* helpers.vhdl:244:32  */
  assign n4821_o = |(n4820_o);
  /* helpers.vhdl:244:28  */
  assign n4822_o = n4819_o | n4821_o;
  /* helpers.vhdl:244:36  */
  assign n4823_o = n4676_o[51:50];
  /* helpers.vhdl:244:32  */
  assign n4824_o = |(n4823_o);
  /* helpers.vhdl:244:28  */
  assign n4825_o = n4822_o | n4824_o;
  /* helpers.vhdl:244:36  */
  assign n4826_o = n4676_o[55:54];
  /* helpers.vhdl:244:32  */
  assign n4827_o = |(n4826_o);
  /* helpers.vhdl:244:28  */
  assign n4828_o = n4825_o | n4827_o;
  /* helpers.vhdl:244:36  */
  assign n4829_o = n4676_o[59:58];
  /* helpers.vhdl:244:32  */
  assign n4830_o = |(n4829_o);
  /* helpers.vhdl:244:28  */
  assign n4831_o = n4828_o | n4830_o;
  /* helpers.vhdl:244:36  */
  assign n4832_o = n4676_o[63:62];
  /* helpers.vhdl:244:32  */
  assign n4833_o = |(n4832_o);
  /* helpers.vhdl:244:28  */
  assign n4834_o = n4831_o | n4833_o;
  /* helpers.vhdl:244:36  */
  assign n4836_o = n4676_o[7:4];
  /* helpers.vhdl:244:32  */
  assign n4837_o = |(n4836_o);
  /* helpers.vhdl:244:28  */
  assign n4839_o = 1'b0 | n4837_o;
  /* helpers.vhdl:244:36  */
  assign n4841_o = n4676_o[15:12];
  /* helpers.vhdl:244:32  */
  assign n4842_o = |(n4841_o);
  /* helpers.vhdl:244:28  */
  assign n4843_o = n4839_o | n4842_o;
  /* helpers.vhdl:244:36  */
  assign n4844_o = n4676_o[23:20];
  /* helpers.vhdl:244:32  */
  assign n4845_o = |(n4844_o);
  /* helpers.vhdl:244:28  */
  assign n4846_o = n4843_o | n4845_o;
  /* helpers.vhdl:244:36  */
  assign n4847_o = n4676_o[31:28];
  /* helpers.vhdl:244:32  */
  assign n4848_o = |(n4847_o);
  /* helpers.vhdl:244:28  */
  assign n4849_o = n4846_o | n4848_o;
  /* helpers.vhdl:244:36  */
  assign n4850_o = n4676_o[39:36];
  /* helpers.vhdl:244:32  */
  assign n4851_o = |(n4850_o);
  /* helpers.vhdl:244:28  */
  assign n4852_o = n4849_o | n4851_o;
  /* helpers.vhdl:244:36  */
  assign n4853_o = n4676_o[47:44];
  /* helpers.vhdl:244:32  */
  assign n4854_o = |(n4853_o);
  /* helpers.vhdl:244:28  */
  assign n4855_o = n4852_o | n4854_o;
  /* helpers.vhdl:244:36  */
  assign n4856_o = n4676_o[55:52];
  /* helpers.vhdl:244:32  */
  assign n4857_o = |(n4856_o);
  /* helpers.vhdl:244:28  */
  assign n4858_o = n4855_o | n4857_o;
  /* helpers.vhdl:244:36  */
  assign n4859_o = n4676_o[63:60];
  /* helpers.vhdl:244:32  */
  assign n4860_o = |(n4859_o);
  /* helpers.vhdl:244:28  */
  assign n4861_o = n4858_o | n4860_o;
  /* helpers.vhdl:244:36  */
  assign n4863_o = n4676_o[15:8];
  /* helpers.vhdl:244:32  */
  assign n4864_o = |(n4863_o);
  /* helpers.vhdl:244:28  */
  assign n4866_o = 1'b0 | n4864_o;
  /* helpers.vhdl:244:36  */
  assign n4868_o = n4676_o[31:24];
  /* helpers.vhdl:244:32  */
  assign n4869_o = |(n4868_o);
  /* helpers.vhdl:244:28  */
  assign n4870_o = n4866_o | n4869_o;
  /* helpers.vhdl:244:36  */
  assign n4871_o = n4676_o[47:40];
  /* helpers.vhdl:244:32  */
  assign n4872_o = |(n4871_o);
  /* helpers.vhdl:244:28  */
  assign n4873_o = n4870_o | n4872_o;
  /* helpers.vhdl:244:36  */
  assign n4874_o = n4676_o[63:56];
  /* helpers.vhdl:244:32  */
  assign n4875_o = |(n4874_o);
  /* helpers.vhdl:244:28  */
  assign n4876_o = n4873_o | n4875_o;
  /* helpers.vhdl:244:36  */
  assign n4878_o = n4676_o[31:16];
  /* helpers.vhdl:244:32  */
  assign n4879_o = |(n4878_o);
  /* helpers.vhdl:244:28  */
  assign n4881_o = 1'b0 | n4879_o;
  /* helpers.vhdl:244:36  */
  assign n4883_o = n4676_o[63:48];
  /* helpers.vhdl:244:32  */
  assign n4884_o = |(n4883_o);
  /* helpers.vhdl:244:28  */
  assign n4885_o = n4881_o | n4884_o;
  /* helpers.vhdl:244:36  */
  assign n4887_o = n4676_o[63:32];
  /* helpers.vhdl:244:32  */
  assign n4888_o = |(n4887_o);
  /* helpers.vhdl:244:28  */
  assign n4890_o = 1'b0 | n4888_o;
  assign n4892_o = {n4890_o, n4885_o, n4876_o, n4861_o, n4834_o, n4782_o};
  /* helpers.vhdl:287:19  */
  assign n4894_o = n4673_o[5:2];
  /* helpers.vhdl:287:38  */
  assign n4895_o = n4892_o[1:0];
  /* helpers.vhdl:287:32  */
  assign n4896_o = {n4894_o, n4895_o};
  /* xics.vhdl:308:17  */
  assign n4899_o = n4896_o[3:0];
  /* xics.vhdl:282:16  */
  assign n4909_o = n4155_o == 3'b111;
  assign n4911_o = n4910_o[7:3];
  assign n4912_o = {n4911_o, n4155_o};
  /* xics.vhdl:282:9  */
  assign n4914_o = n4909_o ? 8'b11111111 : n4912_o;
  /* xics.vhdl:392:9  */
  always @(posedge clk)
    n4918_q <= n3237_o;
  /* xics.vhdl:392:9  */
  assign n4919_o = {n4914_o, n4899_o};
  /* xics.vhdl:350:9  */
  always @(posedge clk)
    n4920_q <= int_level_in;
  /* xics.vhdl:365:9  */
  always @(posedge clk)
    n4921_q <= n3173_o;
  /* xics.vhdl:365:9  */
  assign n4922_o = {1'b0, n4921_q};
  /* xics.vhdl:417:9  */
  always @(posedge clk)
    n4923_q <= icp_out_next;
  /* xics.vhdl:224:9  */
  assign n4924_o = int_level_l[0];
  /* xics.vhdl:221:9  */
  assign n4925_o = int_level_l[1];
  assign n4926_o = int_level_l[2];
  assign n4927_o = int_level_l[3];
  assign n4928_o = int_level_l[4];
  /* xics.vhdl:280:18  */
  assign n4929_o = int_level_l[5];
  assign n4930_o = int_level_l[6];
  /* xics.vhdl:279:14  */
  assign n4931_o = int_level_l[7];
  /* xics.vhdl:279:14  */
  assign n4932_o = int_level_l[8];
  assign n4933_o = int_level_l[9];
  /* xics.vhdl:279:14  */
  assign n4934_o = int_level_l[10];
  /* xics.vhdl:446:20  */
  assign n4935_o = int_level_l[11];
  assign n4936_o = int_level_l[12];
  assign n4937_o = int_level_l[13];
  assign n4938_o = int_level_l[14];
  assign n4939_o = int_level_l[15];
  /* xics.vhdl:369:38  */
  assign n4940_o = reg_idx[1:0];
  /* xics.vhdl:369:38  */
  always @*
    case (n4940_o)
      2'b00: n4941_o = n4924_o;
      2'b01: n4941_o = n4925_o;
      2'b10: n4941_o = n4926_o;
      2'b11: n4941_o = n4927_o;
    endcase
  /* xics.vhdl:369:38  */
  assign n4942_o = reg_idx[1:0];
  /* xics.vhdl:369:38  */
  always @*
    case (n4942_o)
      2'b00: n4943_o = n4928_o;
      2'b01: n4943_o = n4929_o;
      2'b10: n4943_o = n4930_o;
      2'b11: n4943_o = n4931_o;
    endcase
  /* xics.vhdl:369:38  */
  assign n4944_o = reg_idx[1:0];
  /* xics.vhdl:369:38  */
  always @*
    case (n4944_o)
      2'b00: n4945_o = n4932_o;
      2'b01: n4945_o = n4933_o;
      2'b10: n4945_o = n4934_o;
      2'b11: n4945_o = n4935_o;
    endcase
  /* xics.vhdl:369:38  */
  assign n4946_o = reg_idx[1:0];
  /* xics.vhdl:369:38  */
  always @*
    case (n4946_o)
      2'b00: n4947_o = n4936_o;
      2'b01: n4947_o = n4937_o;
      2'b10: n4947_o = n4938_o;
      2'b11: n4947_o = n4939_o;
    endcase
  /* xics.vhdl:369:38  */
  assign n4948_o = reg_idx[3:2];
  /* xics.vhdl:369:38  */
  always @*
    case (n4948_o)
      2'b00: n4949_o = n4941_o;
      2'b01: n4949_o = n4943_o;
      2'b10: n4949_o = n4945_o;
      2'b11: n4949_o = n4947_o;
    endcase
  /* xics.vhdl:369:38  */
  assign n4950_o = int_level_l[0];
  /* xics.vhdl:369:39  */
  assign n4951_o = int_level_l[1];
  assign n4952_o = int_level_l[2];
  assign n4953_o = int_level_l[3];
  /* helpers.vhdl:237:18  */
  assign n4954_o = int_level_l[4];
  assign n4955_o = int_level_l[5];
  /* helpers.vhdl:236:18  */
  assign n4956_o = int_level_l[6];
  assign n4957_o = int_level_l[7];
  /* helpers.vhdl:235:18  */
  assign n4958_o = int_level_l[8];
  assign n4959_o = int_level_l[9];
  /* helpers.vhdl:234:18  */
  assign n4960_o = int_level_l[10];
  assign n4961_o = int_level_l[11];
  /* helpers.vhdl:30:14  */
  assign n4962_o = int_level_l[12];
  /* helpers.vhdl:30:14  */
  assign n4963_o = int_level_l[13];
  assign n4964_o = int_level_l[14];
  /* helpers.vhdl:30:14  */
  assign n4965_o = int_level_l[15];
  /* xics.vhdl:371:38  */
  assign n4966_o = reg_idx[1:0];
  /* xics.vhdl:371:38  */
  always @*
    case (n4966_o)
      2'b00: n4967_o = n4950_o;
      2'b01: n4967_o = n4951_o;
      2'b10: n4967_o = n4952_o;
      2'b11: n4967_o = n4953_o;
    endcase
  /* xics.vhdl:371:38  */
  assign n4968_o = reg_idx[1:0];
  /* xics.vhdl:371:38  */
  always @*
    case (n4968_o)
      2'b00: n4969_o = n4954_o;
      2'b01: n4969_o = n4955_o;
      2'b10: n4969_o = n4956_o;
      2'b11: n4969_o = n4957_o;
    endcase
  /* xics.vhdl:371:38  */
  assign n4970_o = reg_idx[1:0];
  /* xics.vhdl:371:38  */
  always @*
    case (n4970_o)
      2'b00: n4971_o = n4958_o;
      2'b01: n4971_o = n4959_o;
      2'b10: n4971_o = n4960_o;
      2'b11: n4971_o = n4961_o;
    endcase
  /* xics.vhdl:371:38  */
  assign n4972_o = reg_idx[1:0];
  /* xics.vhdl:371:38  */
  always @*
    case (n4972_o)
      2'b00: n4973_o = n4962_o;
      2'b01: n4973_o = n4963_o;
      2'b10: n4973_o = n4964_o;
      2'b11: n4973_o = n4965_o;
    endcase
  /* xics.vhdl:371:38  */
  assign n4974_o = reg_idx[3:2];
  /* xics.vhdl:371:38  */
  always @*
    case (n4974_o)
      2'b00: n4975_o = n4967_o;
      2'b01: n4975_o = n4969_o;
      2'b10: n4975_o = n4971_o;
      2'b11: n4975_o = n4973_o;
    endcase
  /* xics.vhdl:371:38  */
  assign n4976_o = xives[2:0];
  /* xics.vhdl:371:39  */
  assign n4977_o = xives[5:3];
  assign n4978_o = xives[8:6];
  assign n4979_o = xives[11:9];
  assign n4980_o = xives[14:12];
  /* helpers.vhdl:259:18  */
  assign n4981_o = xives[17:15];
  assign n4982_o = xives[20:18];
  /* helpers.vhdl:258:18  */
  assign n4983_o = xives[23:21];
  assign n4984_o = xives[26:24];
  /* helpers.vhdl:257:18  */
  assign n4985_o = xives[29:27];
  assign n4986_o = xives[32:30];
  /* helpers.vhdl:256:18  */
  assign n4987_o = xives[35:33];
  assign n4988_o = xives[38:36];
  /* helpers.vhdl:31:14  */
  assign n4989_o = xives[41:39];
  /* helpers.vhdl:31:14  */
  assign n4990_o = xives[44:42];
  assign n4991_o = xives[47:45];
  /* xics.vhdl:374:44  */
  assign n4992_o = n3128_o[1:0];
  /* xics.vhdl:374:44  */
  always @*
    case (n4992_o)
      2'b00: n4993_o = n4976_o;
      2'b01: n4993_o = n4977_o;
      2'b10: n4993_o = n4978_o;
      2'b11: n4993_o = n4979_o;
    endcase
  /* xics.vhdl:374:44  */
  assign n4994_o = n3128_o[1:0];
  /* xics.vhdl:374:44  */
  always @*
    case (n4994_o)
      2'b00: n4995_o = n4980_o;
      2'b01: n4995_o = n4981_o;
      2'b10: n4995_o = n4982_o;
      2'b11: n4995_o = n4983_o;
    endcase
  /* xics.vhdl:374:44  */
  assign n4996_o = n3128_o[1:0];
  /* xics.vhdl:374:44  */
  always @*
    case (n4996_o)
      2'b00: n4997_o = n4984_o;
      2'b01: n4997_o = n4985_o;
      2'b10: n4997_o = n4986_o;
      2'b11: n4997_o = n4987_o;
    endcase
  /* xics.vhdl:374:44  */
  assign n4998_o = n3128_o[1:0];
  /* xics.vhdl:374:44  */
  always @*
    case (n4998_o)
      2'b00: n4999_o = n4988_o;
      2'b01: n4999_o = n4989_o;
      2'b10: n4999_o = n4990_o;
      2'b11: n4999_o = n4991_o;
    endcase
  /* xics.vhdl:374:44  */
  assign n5000_o = n3128_o[3:2];
  /* xics.vhdl:374:44  */
  always @*
    case (n5000_o)
      2'b00: n5001_o = n4993_o;
      2'b01: n5001_o = n4995_o;
      2'b10: n5001_o = n4997_o;
      2'b11: n5001_o = n4999_o;
    endcase
  /* xics.vhdl:401:21  */
  assign n5002_o = n3216_o[3];
  /* xics.vhdl:401:21  */
  assign n5003_o = ~n5002_o;
  /* xics.vhdl:401:21  */
  assign n5004_o = n3216_o[2];
  /* xics.vhdl:401:21  */
  assign n5005_o = ~n5004_o;
  /* xics.vhdl:401:21  */
  assign n5006_o = n5003_o & n5005_o;
  /* xics.vhdl:401:21  */
  assign n5007_o = n5003_o & n5004_o;
  /* xics.vhdl:401:21  */
  assign n5008_o = n5002_o & n5005_o;
  /* xics.vhdl:401:21  */
  assign n5009_o = n5002_o & n5004_o;
  /* xics.vhdl:401:21  */
  assign n5010_o = n3216_o[1];
  /* xics.vhdl:401:21  */
  assign n5011_o = ~n5010_o;
  /* xics.vhdl:401:21  */
  assign n5012_o = n5006_o & n5011_o;
  /* xics.vhdl:401:21  */
  assign n5013_o = n5006_o & n5010_o;
  /* xics.vhdl:401:21  */
  assign n5014_o = n5007_o & n5011_o;
  /* xics.vhdl:401:21  */
  assign n5015_o = n5007_o & n5010_o;
  /* xics.vhdl:401:21  */
  assign n5016_o = n5008_o & n5011_o;
  /* xics.vhdl:401:21  */
  assign n5017_o = n5008_o & n5010_o;
  /* xics.vhdl:401:21  */
  assign n5018_o = n5009_o & n5011_o;
  /* xics.vhdl:401:21  */
  assign n5019_o = n5009_o & n5010_o;
  /* xics.vhdl:401:21  */
  assign n5020_o = n3216_o[0];
  /* xics.vhdl:401:21  */
  assign n5021_o = ~n5020_o;
  /* xics.vhdl:401:21  */
  assign n5022_o = n5012_o & n5021_o;
  /* xics.vhdl:401:21  */
  assign n5023_o = n5012_o & n5020_o;
  /* xics.vhdl:401:21  */
  assign n5024_o = n5013_o & n5021_o;
  /* xics.vhdl:401:21  */
  assign n5025_o = n5013_o & n5020_o;
  /* xics.vhdl:401:21  */
  assign n5026_o = n5014_o & n5021_o;
  /* xics.vhdl:401:21  */
  assign n5027_o = n5014_o & n5020_o;
  /* xics.vhdl:401:21  */
  assign n5028_o = n5015_o & n5021_o;
  /* xics.vhdl:401:21  */
  assign n5029_o = n5015_o & n5020_o;
  /* xics.vhdl:401:21  */
  assign n5030_o = n5016_o & n5021_o;
  /* xics.vhdl:401:21  */
  assign n5031_o = n5016_o & n5020_o;
  /* xics.vhdl:401:21  */
  assign n5032_o = n5017_o & n5021_o;
  /* xics.vhdl:401:21  */
  assign n5033_o = n5017_o & n5020_o;
  /* xics.vhdl:401:21  */
  assign n5034_o = n5018_o & n5021_o;
  /* xics.vhdl:401:21  */
  assign n5035_o = n5018_o & n5020_o;
  /* xics.vhdl:401:21  */
  assign n5036_o = n5019_o & n5021_o;
  /* xics.vhdl:401:21  */
  assign n5037_o = n5019_o & n5020_o;
  assign n5038_o = xives[2:0];
  /* xics.vhdl:401:21  */
  assign n5039_o = n5022_o ? n3232_o : n5038_o;
  assign n5040_o = xives[5:3];
  /* xics.vhdl:401:21  */
  assign n5041_o = n5023_o ? n3232_o : n5040_o;
  assign n5042_o = xives[8:6];
  /* xics.vhdl:401:21  */
  assign n5043_o = n5024_o ? n3232_o : n5042_o;
  assign n5044_o = xives[11:9];
  /* xics.vhdl:401:21  */
  assign n5045_o = n5025_o ? n3232_o : n5044_o;
  assign n5046_o = xives[14:12];
  /* xics.vhdl:401:21  */
  assign n5047_o = n5026_o ? n3232_o : n5046_o;
  assign n5048_o = xives[17:15];
  /* xics.vhdl:401:21  */
  assign n5049_o = n5027_o ? n3232_o : n5048_o;
  assign n5050_o = xives[20:18];
  /* xics.vhdl:401:21  */
  assign n5051_o = n5028_o ? n3232_o : n5050_o;
  /* helpers.vhdl:237:18  */
  assign n5052_o = xives[23:21];
  /* xics.vhdl:401:21  */
  assign n5053_o = n5029_o ? n3232_o : n5052_o;
  /* helpers.vhdl:236:18  */
  assign n5054_o = xives[26:24];
  /* xics.vhdl:401:21  */
  assign n5055_o = n5030_o ? n3232_o : n5054_o;
  /* helpers.vhdl:235:18  */
  assign n5056_o = xives[29:27];
  /* xics.vhdl:401:21  */
  assign n5057_o = n5031_o ? n3232_o : n5056_o;
  /* helpers.vhdl:234:18  */
  assign n5058_o = xives[32:30];
  /* xics.vhdl:401:21  */
  assign n5059_o = n5032_o ? n3232_o : n5058_o;
  /* helpers.vhdl:30:14  */
  assign n5060_o = xives[35:33];
  /* xics.vhdl:401:21  */
  assign n5061_o = n5033_o ? n3232_o : n5060_o;
  assign n5062_o = xives[38:36];
  /* xics.vhdl:401:21  */
  assign n5063_o = n5034_o ? n3232_o : n5062_o;
  assign n5064_o = xives[41:39];
  /* xics.vhdl:401:21  */
  assign n5065_o = n5035_o ? n3232_o : n5064_o;
  assign n5066_o = xives[44:42];
  /* xics.vhdl:401:21  */
  assign n5067_o = n5036_o ? n3232_o : n5066_o;
  assign n5068_o = xives[47:45];
  /* xics.vhdl:401:21  */
  assign n5069_o = n5037_o ? n3232_o : n5068_o;
  assign n5070_o = {n5069_o, n5067_o, n5065_o, n5063_o, n5061_o, n5059_o, n5057_o, n5055_o, n5053_o, n5051_o, n5049_o, n5047_o, n5045_o, n5043_o, n5041_o, n5039_o};
  /* xics.vhdl:295:9  */
  assign n5071_o = n3252_o[2];
  /* xics.vhdl:295:9  */
  assign n5072_o = ~n5071_o;
  /* xics.vhdl:295:9  */
  assign n5073_o = n3252_o[1];
  /* xics.vhdl:295:9  */
  assign n5074_o = ~n5073_o;
  /* xics.vhdl:295:9  */
  assign n5075_o = n5072_o & n5074_o;
  /* xics.vhdl:295:9  */
  assign n5076_o = n5072_o & n5073_o;
  /* xics.vhdl:295:9  */
  assign n5077_o = n5071_o & n5074_o;
  /* xics.vhdl:295:9  */
  assign n5078_o = n5071_o & n5073_o;
  /* xics.vhdl:295:9  */
  assign n5079_o = n3252_o[0];
  /* xics.vhdl:295:9  */
  assign n5080_o = ~n5079_o;
  /* xics.vhdl:295:9  */
  assign n5081_o = n5075_o & n5080_o;
  /* xics.vhdl:295:9  */
  assign n5082_o = n5075_o & n5079_o;
  /* xics.vhdl:295:9  */
  assign n5083_o = n5076_o & n5080_o;
  /* xics.vhdl:295:9  */
  assign n5084_o = n5076_o & n5079_o;
  /* xics.vhdl:295:9  */
  assign n5085_o = n5077_o & n5080_o;
  /* xics.vhdl:295:9  */
  assign n5086_o = n5077_o & n5079_o;
  /* xics.vhdl:295:9  */
  assign n5087_o = n5078_o & n5080_o;
  /* xics.vhdl:295:9  */
  assign n5088_o = n5078_o & n5079_o;
  assign n5089_o = n3260_o[0];
  /* xics.vhdl:295:9  */
  assign n5090_o = n5081_o ? 1'b1 : n5089_o;
  assign n5091_o = n3260_o[1];
  /* xics.vhdl:295:9  */
  assign n5092_o = n5082_o ? 1'b1 : n5091_o;
  assign n5093_o = n3260_o[2];
  /* xics.vhdl:295:9  */
  assign n5094_o = n5083_o ? 1'b1 : n5093_o;
  assign n5095_o = n3260_o[3];
  /* xics.vhdl:295:9  */
  assign n5096_o = n5084_o ? 1'b1 : n5095_o;
  assign n5097_o = n3260_o[4];
  /* xics.vhdl:295:9  */
  assign n5098_o = n5085_o ? 1'b1 : n5097_o;
  assign n5099_o = n3260_o[5];
  /* xics.vhdl:295:9  */
  assign n5100_o = n5086_o ? 1'b1 : n5099_o;
  assign n5101_o = n3260_o[6];
  /* xics.vhdl:295:9  */
  assign n5102_o = n5087_o ? 1'b1 : n5101_o;
  assign n5103_o = n3260_o[7];
  /* xics.vhdl:295:9  */
  assign n5104_o = n5088_o ? 1'b1 : n5103_o;
  assign n5105_o = {n5104_o, n5102_o, n5100_o, n5098_o, n5096_o, n5094_o, n5092_o, n5090_o};
  /* xics.vhdl:295:9  */
  assign n5106_o = n3272_o[2];
  /* xics.vhdl:295:9  */
  assign n5107_o = ~n5106_o;
  /* xics.vhdl:295:9  */
  assign n5108_o = n3272_o[1];
  /* xics.vhdl:295:9  */
  assign n5109_o = ~n5108_o;
  /* xics.vhdl:295:9  */
  assign n5110_o = n5107_o & n5109_o;
  /* xics.vhdl:295:9  */
  assign n5111_o = n5107_o & n5108_o;
  /* xics.vhdl:295:9  */
  assign n5112_o = n5106_o & n5109_o;
  /* xics.vhdl:295:9  */
  assign n5113_o = n5106_o & n5108_o;
  /* xics.vhdl:295:9  */
  assign n5114_o = n3272_o[0];
  /* xics.vhdl:295:9  */
  assign n5115_o = ~n5114_o;
  /* xics.vhdl:295:9  */
  assign n5116_o = n5110_o & n5115_o;
  /* xics.vhdl:295:9  */
  assign n5117_o = n5110_o & n5114_o;
  /* xics.vhdl:295:9  */
  assign n5118_o = n5111_o & n5115_o;
  /* xics.vhdl:295:9  */
  assign n5119_o = n5111_o & n5114_o;
  /* xics.vhdl:295:9  */
  assign n5120_o = n5112_o & n5115_o;
  /* xics.vhdl:295:9  */
  assign n5121_o = n5112_o & n5114_o;
  /* xics.vhdl:295:9  */
  assign n5122_o = n5113_o & n5115_o;
  /* xics.vhdl:295:9  */
  assign n5123_o = n5113_o & n5114_o;
  /* xics.vhdl:292:18  */
  assign n5124_o = n3280_o[0];
  /* xics.vhdl:295:9  */
  assign n5125_o = n5116_o ? 1'b1 : n5124_o;
  /* xics.vhdl:291:14  */
  assign n5126_o = n3280_o[1];
  /* xics.vhdl:295:9  */
  assign n5127_o = n5117_o ? 1'b1 : n5126_o;
  assign n5128_o = n3280_o[2];
  /* xics.vhdl:295:9  */
  assign n5129_o = n5118_o ? 1'b1 : n5128_o;
  assign n5130_o = n3280_o[3];
  /* xics.vhdl:295:9  */
  assign n5131_o = n5119_o ? 1'b1 : n5130_o;
  /* xics.vhdl:292:18  */
  assign n5132_o = n3280_o[4];
  /* xics.vhdl:295:9  */
  assign n5133_o = n5120_o ? 1'b1 : n5132_o;
  /* xics.vhdl:291:14  */
  assign n5134_o = n3280_o[5];
  /* xics.vhdl:295:9  */
  assign n5135_o = n5121_o ? 1'b1 : n5134_o;
  assign n5136_o = n3280_o[6];
  /* xics.vhdl:295:9  */
  assign n5137_o = n5122_o ? 1'b1 : n5136_o;
  assign n5138_o = n3280_o[7];
  /* xics.vhdl:295:9  */
  assign n5139_o = n5123_o ? 1'b1 : n5138_o;
  /* xics.vhdl:292:18  */
  assign n5140_o = {n5139_o, n5137_o, n5135_o, n5133_o, n5131_o, n5129_o, n5127_o, n5125_o};
  /* xics.vhdl:295:9  */
  assign n5141_o = n3289_o[2];
  /* xics.vhdl:295:9  */
  assign n5142_o = ~n5141_o;
  /* xics.vhdl:295:9  */
  assign n5143_o = n3289_o[1];
  /* xics.vhdl:295:9  */
  assign n5144_o = ~n5143_o;
  /* xics.vhdl:295:9  */
  assign n5145_o = n5142_o & n5144_o;
  /* xics.vhdl:295:9  */
  assign n5146_o = n5142_o & n5143_o;
  /* xics.vhdl:295:9  */
  assign n5147_o = n5141_o & n5144_o;
  /* xics.vhdl:295:9  */
  assign n5148_o = n5141_o & n5143_o;
  /* xics.vhdl:295:9  */
  assign n5149_o = n3289_o[0];
  /* xics.vhdl:295:9  */
  assign n5150_o = ~n5149_o;
  /* xics.vhdl:295:9  */
  assign n5151_o = n5145_o & n5150_o;
  /* xics.vhdl:295:9  */
  assign n5152_o = n5145_o & n5149_o;
  /* xics.vhdl:295:9  */
  assign n5153_o = n5146_o & n5150_o;
  /* xics.vhdl:295:9  */
  assign n5154_o = n5146_o & n5149_o;
  /* xics.vhdl:295:9  */
  assign n5155_o = n5147_o & n5150_o;
  /* xics.vhdl:295:9  */
  assign n5156_o = n5147_o & n5149_o;
  /* xics.vhdl:295:9  */
  assign n5157_o = n5148_o & n5150_o;
  /* xics.vhdl:295:9  */
  assign n5158_o = n5148_o & n5149_o;
  assign n5159_o = n3297_o[0];
  /* xics.vhdl:295:9  */
  assign n5160_o = n5151_o ? 1'b1 : n5159_o;
  /* xics.vhdl:291:14  */
  assign n5161_o = n3297_o[1];
  /* xics.vhdl:295:9  */
  assign n5162_o = n5152_o ? 1'b1 : n5161_o;
  /* xics.vhdl:291:14  */
  assign n5163_o = n3297_o[2];
  /* xics.vhdl:295:9  */
  assign n5164_o = n5153_o ? 1'b1 : n5163_o;
  /* xics.vhdl:295:11  */
  assign n5165_o = n3297_o[3];
  /* xics.vhdl:295:9  */
  assign n5166_o = n5154_o ? 1'b1 : n5165_o;
  assign n5167_o = n3297_o[4];
  /* xics.vhdl:295:9  */
  assign n5168_o = n5155_o ? 1'b1 : n5167_o;
  /* xics.vhdl:291:14  */
  assign n5169_o = n3297_o[5];
  /* xics.vhdl:295:9  */
  assign n5170_o = n5156_o ? 1'b1 : n5169_o;
  /* xics.vhdl:291:14  */
  assign n5171_o = n3297_o[6];
  /* xics.vhdl:295:9  */
  assign n5172_o = n5157_o ? 1'b1 : n5171_o;
  /* xics.vhdl:295:11  */
  assign n5173_o = n3297_o[7];
  /* xics.vhdl:295:9  */
  assign n5174_o = n5158_o ? 1'b1 : n5173_o;
  assign n5175_o = {n5174_o, n5172_o, n5170_o, n5168_o, n5166_o, n5164_o, n5162_o, n5160_o};
  /* xics.vhdl:295:9  */
  assign n5176_o = n3306_o[2];
  /* xics.vhdl:295:9  */
  assign n5177_o = ~n5176_o;
  /* xics.vhdl:295:9  */
  assign n5178_o = n3306_o[1];
  /* xics.vhdl:295:9  */
  assign n5179_o = ~n5178_o;
  /* xics.vhdl:295:9  */
  assign n5180_o = n5177_o & n5179_o;
  /* xics.vhdl:295:9  */
  assign n5181_o = n5177_o & n5178_o;
  /* xics.vhdl:295:9  */
  assign n5182_o = n5176_o & n5179_o;
  /* xics.vhdl:295:9  */
  assign n5183_o = n5176_o & n5178_o;
  /* xics.vhdl:295:9  */
  assign n5184_o = n3306_o[0];
  /* xics.vhdl:295:9  */
  assign n5185_o = ~n5184_o;
  /* xics.vhdl:295:9  */
  assign n5186_o = n5180_o & n5185_o;
  /* xics.vhdl:295:9  */
  assign n5187_o = n5180_o & n5184_o;
  /* xics.vhdl:295:9  */
  assign n5188_o = n5181_o & n5185_o;
  /* xics.vhdl:295:9  */
  assign n5189_o = n5181_o & n5184_o;
  /* xics.vhdl:295:9  */
  assign n5190_o = n5182_o & n5185_o;
  /* xics.vhdl:295:9  */
  assign n5191_o = n5182_o & n5184_o;
  /* xics.vhdl:295:9  */
  assign n5192_o = n5183_o & n5185_o;
  /* xics.vhdl:295:9  */
  assign n5193_o = n5183_o & n5184_o;
  /* xics.vhdl:291:14  */
  assign n5194_o = n3314_o[0];
  /* xics.vhdl:295:9  */
  assign n5195_o = n5186_o ? 1'b1 : n5194_o;
  assign n5196_o = n3314_o[1];
  /* xics.vhdl:295:9  */
  assign n5197_o = n5187_o ? 1'b1 : n5196_o;
  assign n5198_o = n3314_o[2];
  /* xics.vhdl:295:9  */
  assign n5199_o = n5188_o ? 1'b1 : n5198_o;
  /* xics.vhdl:292:18  */
  assign n5200_o = n3314_o[3];
  /* xics.vhdl:295:9  */
  assign n5201_o = n5189_o ? 1'b1 : n5200_o;
  /* xics.vhdl:291:14  */
  assign n5202_o = n3314_o[4];
  /* xics.vhdl:295:9  */
  assign n5203_o = n5190_o ? 1'b1 : n5202_o;
  assign n5204_o = n3314_o[5];
  /* xics.vhdl:295:9  */
  assign n5205_o = n5191_o ? 1'b1 : n5204_o;
  assign n5206_o = n3314_o[6];
  /* xics.vhdl:295:9  */
  assign n5207_o = n5192_o ? 1'b1 : n5206_o;
  /* xics.vhdl:292:18  */
  assign n5208_o = n3314_o[7];
  /* xics.vhdl:295:9  */
  assign n5209_o = n5193_o ? 1'b1 : n5208_o;
  /* xics.vhdl:291:14  */
  assign n5210_o = {n5209_o, n5207_o, n5205_o, n5203_o, n5201_o, n5199_o, n5197_o, n5195_o};
  /* xics.vhdl:295:9  */
  assign n5211_o = n3323_o[2];
  /* xics.vhdl:295:9  */
  assign n5212_o = ~n5211_o;
  /* xics.vhdl:295:9  */
  assign n5213_o = n3323_o[1];
  /* xics.vhdl:295:9  */
  assign n5214_o = ~n5213_o;
  /* xics.vhdl:295:9  */
  assign n5215_o = n5212_o & n5214_o;
  /* xics.vhdl:295:9  */
  assign n5216_o = n5212_o & n5213_o;
  /* xics.vhdl:295:9  */
  assign n5217_o = n5211_o & n5214_o;
  /* xics.vhdl:295:9  */
  assign n5218_o = n5211_o & n5213_o;
  /* xics.vhdl:295:9  */
  assign n5219_o = n3323_o[0];
  /* xics.vhdl:295:9  */
  assign n5220_o = ~n5219_o;
  /* xics.vhdl:295:9  */
  assign n5221_o = n5215_o & n5220_o;
  /* xics.vhdl:295:9  */
  assign n5222_o = n5215_o & n5219_o;
  /* xics.vhdl:295:9  */
  assign n5223_o = n5216_o & n5220_o;
  /* xics.vhdl:295:9  */
  assign n5224_o = n5216_o & n5219_o;
  /* xics.vhdl:295:9  */
  assign n5225_o = n5217_o & n5220_o;
  /* xics.vhdl:295:9  */
  assign n5226_o = n5217_o & n5219_o;
  /* xics.vhdl:295:9  */
  assign n5227_o = n5218_o & n5220_o;
  /* xics.vhdl:295:9  */
  assign n5228_o = n5218_o & n5219_o;
  /* xics.vhdl:291:14  */
  assign n5229_o = n3331_o[0];
  /* xics.vhdl:295:9  */
  assign n5230_o = n5221_o ? 1'b1 : n5229_o;
  /* xics.vhdl:291:14  */
  assign n5231_o = n3331_o[1];
  /* xics.vhdl:295:9  */
  assign n5232_o = n5222_o ? 1'b1 : n5231_o;
  /* xics.vhdl:295:11  */
  assign n5233_o = n3331_o[2];
  /* xics.vhdl:295:9  */
  assign n5234_o = n5223_o ? 1'b1 : n5233_o;
  assign n5235_o = n3331_o[3];
  /* xics.vhdl:295:9  */
  assign n5236_o = n5224_o ? 1'b1 : n5235_o;
  /* xics.vhdl:291:14  */
  assign n5237_o = n3331_o[4];
  /* xics.vhdl:295:9  */
  assign n5238_o = n5225_o ? 1'b1 : n5237_o;
  /* xics.vhdl:291:14  */
  assign n5239_o = n3331_o[5];
  /* xics.vhdl:295:9  */
  assign n5240_o = n5226_o ? 1'b1 : n5239_o;
  /* xics.vhdl:295:11  */
  assign n5241_o = n3331_o[6];
  /* xics.vhdl:295:9  */
  assign n5242_o = n5227_o ? 1'b1 : n5241_o;
  assign n5243_o = n3331_o[7];
  /* xics.vhdl:295:9  */
  assign n5244_o = n5228_o ? 1'b1 : n5243_o;
  /* xics.vhdl:291:14  */
  assign n5245_o = {n5244_o, n5242_o, n5240_o, n5238_o, n5236_o, n5234_o, n5232_o, n5230_o};
  /* xics.vhdl:295:9  */
  assign n5246_o = n3340_o[2];
  /* xics.vhdl:295:9  */
  assign n5247_o = ~n5246_o;
  /* xics.vhdl:295:9  */
  assign n5248_o = n3340_o[1];
  /* xics.vhdl:295:9  */
  assign n5249_o = ~n5248_o;
  /* xics.vhdl:295:9  */
  assign n5250_o = n5247_o & n5249_o;
  /* xics.vhdl:295:9  */
  assign n5251_o = n5247_o & n5248_o;
  /* xics.vhdl:295:9  */
  assign n5252_o = n5246_o & n5249_o;
  /* xics.vhdl:295:9  */
  assign n5253_o = n5246_o & n5248_o;
  /* xics.vhdl:295:9  */
  assign n5254_o = n3340_o[0];
  /* xics.vhdl:295:9  */
  assign n5255_o = ~n5254_o;
  /* xics.vhdl:295:9  */
  assign n5256_o = n5250_o & n5255_o;
  /* xics.vhdl:295:9  */
  assign n5257_o = n5250_o & n5254_o;
  /* xics.vhdl:295:9  */
  assign n5258_o = n5251_o & n5255_o;
  /* xics.vhdl:295:9  */
  assign n5259_o = n5251_o & n5254_o;
  /* xics.vhdl:295:9  */
  assign n5260_o = n5252_o & n5255_o;
  /* xics.vhdl:295:9  */
  assign n5261_o = n5252_o & n5254_o;
  /* xics.vhdl:295:9  */
  assign n5262_o = n5253_o & n5255_o;
  /* xics.vhdl:295:9  */
  assign n5263_o = n5253_o & n5254_o;
  /* xics.vhdl:424:18  */
  assign n5264_o = n3348_o[0];
  /* xics.vhdl:295:9  */
  assign n5265_o = n5256_o ? 1'b1 : n5264_o;
  /* xics.vhdl:423:18  */
  assign n5266_o = n3348_o[1];
  /* xics.vhdl:295:9  */
  assign n5267_o = n5257_o ? 1'b1 : n5266_o;
  assign n5268_o = n3348_o[2];
  /* xics.vhdl:295:9  */
  assign n5269_o = n5258_o ? 1'b1 : n5268_o;
  assign n5270_o = n3348_o[3];
  /* xics.vhdl:295:9  */
  assign n5271_o = n5259_o ? 1'b1 : n5270_o;
  assign n5272_o = n3348_o[4];
  /* xics.vhdl:295:9  */
  assign n5273_o = n5260_o ? 1'b1 : n5272_o;
  /* xics.vhdl:267:14  */
  assign n5274_o = n3348_o[5];
  /* xics.vhdl:295:9  */
  assign n5275_o = n5261_o ? 1'b1 : n5274_o;
  /* xics.vhdl:267:14  */
  assign n5276_o = n3348_o[6];
  /* xics.vhdl:295:9  */
  assign n5277_o = n5262_o ? 1'b1 : n5276_o;
  assign n5278_o = n3348_o[7];
  /* xics.vhdl:295:9  */
  assign n5279_o = n5263_o ? 1'b1 : n5278_o;
  assign n5280_o = {n5279_o, n5277_o, n5275_o, n5273_o, n5271_o, n5269_o, n5267_o, n5265_o};
  /* xics.vhdl:295:9  */
  assign n5281_o = n3357_o[2];
  /* xics.vhdl:295:9  */
  assign n5282_o = ~n5281_o;
  /* xics.vhdl:295:9  */
  assign n5283_o = n3357_o[1];
  /* xics.vhdl:295:9  */
  assign n5284_o = ~n5283_o;
  /* xics.vhdl:295:9  */
  assign n5285_o = n5282_o & n5284_o;
  /* xics.vhdl:295:9  */
  assign n5286_o = n5282_o & n5283_o;
  /* xics.vhdl:295:9  */
  assign n5287_o = n5281_o & n5284_o;
  /* xics.vhdl:295:9  */
  assign n5288_o = n5281_o & n5283_o;
  /* xics.vhdl:295:9  */
  assign n5289_o = n3357_o[0];
  /* xics.vhdl:295:9  */
  assign n5290_o = ~n5289_o;
  /* xics.vhdl:295:9  */
  assign n5291_o = n5285_o & n5290_o;
  /* xics.vhdl:295:9  */
  assign n5292_o = n5285_o & n5289_o;
  /* xics.vhdl:295:9  */
  assign n5293_o = n5286_o & n5290_o;
  /* xics.vhdl:295:9  */
  assign n5294_o = n5286_o & n5289_o;
  /* xics.vhdl:295:9  */
  assign n5295_o = n5287_o & n5290_o;
  /* xics.vhdl:295:9  */
  assign n5296_o = n5287_o & n5289_o;
  /* xics.vhdl:295:9  */
  assign n5297_o = n5288_o & n5290_o;
  /* xics.vhdl:295:9  */
  assign n5298_o = n5288_o & n5289_o;
  /* xics.vhdl:249:18  */
  assign n5299_o = n3365_o[0];
  /* xics.vhdl:295:9  */
  assign n5300_o = n5291_o ? 1'b1 : n5299_o;
  /* xics.vhdl:248:14  */
  assign n5301_o = n3365_o[1];
  /* xics.vhdl:295:9  */
  assign n5302_o = n5292_o ? 1'b1 : n5301_o;
  assign n5303_o = n3365_o[2];
  /* xics.vhdl:295:9  */
  assign n5304_o = n5293_o ? 1'b1 : n5303_o;
  assign n5305_o = n3365_o[3];
  /* xics.vhdl:295:9  */
  assign n5306_o = n5294_o ? 1'b1 : n5305_o;
  /* xics.vhdl:280:18  */
  assign n5307_o = n3365_o[4];
  /* xics.vhdl:295:9  */
  assign n5308_o = n5295_o ? 1'b1 : n5307_o;
  /* xics.vhdl:279:14  */
  assign n5309_o = n3365_o[5];
  /* xics.vhdl:295:9  */
  assign n5310_o = n5296_o ? 1'b1 : n5309_o;
  /* xics.vhdl:65:5  */
  assign n5311_o = n3365_o[6];
  /* xics.vhdl:295:9  */
  assign n5312_o = n5297_o ? 1'b1 : n5311_o;
  /* xics.vhdl:362:5  */
  assign n5313_o = n3365_o[7];
  /* xics.vhdl:295:9  */
  assign n5314_o = n5298_o ? 1'b1 : n5313_o;
  assign n5315_o = {n5314_o, n5312_o, n5310_o, n5308_o, n5306_o, n5304_o, n5302_o, n5300_o};
  /* xics.vhdl:295:9  */
  assign n5316_o = n3374_o[2];
  /* xics.vhdl:295:9  */
  assign n5317_o = ~n5316_o;
  /* xics.vhdl:295:9  */
  assign n5318_o = n3374_o[1];
  /* xics.vhdl:295:9  */
  assign n5319_o = ~n5318_o;
  /* xics.vhdl:295:9  */
  assign n5320_o = n5317_o & n5319_o;
  /* xics.vhdl:295:9  */
  assign n5321_o = n5317_o & n5318_o;
  /* xics.vhdl:295:9  */
  assign n5322_o = n5316_o & n5319_o;
  /* xics.vhdl:295:9  */
  assign n5323_o = n5316_o & n5318_o;
  /* xics.vhdl:295:9  */
  assign n5324_o = n3374_o[0];
  /* xics.vhdl:295:9  */
  assign n5325_o = ~n5324_o;
  /* xics.vhdl:295:9  */
  assign n5326_o = n5320_o & n5325_o;
  /* xics.vhdl:295:9  */
  assign n5327_o = n5320_o & n5324_o;
  /* xics.vhdl:295:9  */
  assign n5328_o = n5321_o & n5325_o;
  /* xics.vhdl:295:9  */
  assign n5329_o = n5321_o & n5324_o;
  /* xics.vhdl:295:9  */
  assign n5330_o = n5322_o & n5325_o;
  /* xics.vhdl:295:9  */
  assign n5331_o = n5322_o & n5324_o;
  /* xics.vhdl:295:9  */
  assign n5332_o = n5323_o & n5325_o;
  /* xics.vhdl:295:9  */
  assign n5333_o = n5323_o & n5324_o;
  assign n5334_o = n3382_o[0];
  /* xics.vhdl:295:9  */
  assign n5335_o = n5326_o ? 1'b1 : n5334_o;
  assign n5336_o = n3382_o[1];
  /* xics.vhdl:295:9  */
  assign n5337_o = n5327_o ? 1'b1 : n5336_o;
  assign n5338_o = n3382_o[2];
  /* xics.vhdl:295:9  */
  assign n5339_o = n5328_o ? 1'b1 : n5338_o;
  assign n5340_o = n3382_o[3];
  /* xics.vhdl:295:9  */
  assign n5341_o = n5329_o ? 1'b1 : n5340_o;
  assign n5342_o = n3382_o[4];
  /* xics.vhdl:295:9  */
  assign n5343_o = n5330_o ? 1'b1 : n5342_o;
  assign n5344_o = n3382_o[5];
  /* xics.vhdl:295:9  */
  assign n5345_o = n5331_o ? 1'b1 : n5344_o;
  assign n5346_o = n3382_o[6];
  /* xics.vhdl:295:9  */
  assign n5347_o = n5332_o ? 1'b1 : n5346_o;
  assign n5348_o = n3382_o[7];
  /* xics.vhdl:295:9  */
  assign n5349_o = n5333_o ? 1'b1 : n5348_o;
  assign n5350_o = {n5349_o, n5347_o, n5345_o, n5343_o, n5341_o, n5339_o, n5337_o, n5335_o};
  /* xics.vhdl:295:9  */
  assign n5351_o = n3391_o[2];
  /* xics.vhdl:295:9  */
  assign n5352_o = ~n5351_o;
  /* xics.vhdl:295:9  */
  assign n5353_o = n3391_o[1];
  /* xics.vhdl:295:9  */
  assign n5354_o = ~n5353_o;
  /* xics.vhdl:295:9  */
  assign n5355_o = n5352_o & n5354_o;
  /* xics.vhdl:295:9  */
  assign n5356_o = n5352_o & n5353_o;
  /* xics.vhdl:295:9  */
  assign n5357_o = n5351_o & n5354_o;
  /* xics.vhdl:295:9  */
  assign n5358_o = n5351_o & n5353_o;
  /* xics.vhdl:295:9  */
  assign n5359_o = n3391_o[0];
  /* xics.vhdl:295:9  */
  assign n5360_o = ~n5359_o;
  /* xics.vhdl:295:9  */
  assign n5361_o = n5355_o & n5360_o;
  /* xics.vhdl:295:9  */
  assign n5362_o = n5355_o & n5359_o;
  /* xics.vhdl:295:9  */
  assign n5363_o = n5356_o & n5360_o;
  /* xics.vhdl:295:9  */
  assign n5364_o = n5356_o & n5359_o;
  /* xics.vhdl:295:9  */
  assign n5365_o = n5357_o & n5360_o;
  /* xics.vhdl:295:9  */
  assign n5366_o = n5357_o & n5359_o;
  /* xics.vhdl:295:9  */
  assign n5367_o = n5358_o & n5360_o;
  /* xics.vhdl:295:9  */
  assign n5368_o = n5358_o & n5359_o;
  assign n5369_o = n3399_o[0];
  /* xics.vhdl:295:9  */
  assign n5370_o = n5361_o ? 1'b1 : n5369_o;
  assign n5371_o = n3399_o[1];
  /* xics.vhdl:295:9  */
  assign n5372_o = n5362_o ? 1'b1 : n5371_o;
  assign n5373_o = n3399_o[2];
  /* xics.vhdl:295:9  */
  assign n5374_o = n5363_o ? 1'b1 : n5373_o;
  assign n5375_o = n3399_o[3];
  /* xics.vhdl:295:9  */
  assign n5376_o = n5364_o ? 1'b1 : n5375_o;
  assign n5377_o = n3399_o[4];
  /* xics.vhdl:295:9  */
  assign n5378_o = n5365_o ? 1'b1 : n5377_o;
  assign n5379_o = n3399_o[5];
  /* xics.vhdl:295:9  */
  assign n5380_o = n5366_o ? 1'b1 : n5379_o;
  assign n5381_o = n3399_o[6];
  /* xics.vhdl:295:9  */
  assign n5382_o = n5367_o ? 1'b1 : n5381_o;
  assign n5383_o = n3399_o[7];
  /* xics.vhdl:295:9  */
  assign n5384_o = n5368_o ? 1'b1 : n5383_o;
  assign n5385_o = {n5384_o, n5382_o, n5380_o, n5378_o, n5376_o, n5374_o, n5372_o, n5370_o};
  /* xics.vhdl:295:9  */
  assign n5386_o = n3408_o[2];
  /* xics.vhdl:295:9  */
  assign n5387_o = ~n5386_o;
  /* xics.vhdl:295:9  */
  assign n5388_o = n3408_o[1];
  /* xics.vhdl:295:9  */
  assign n5389_o = ~n5388_o;
  /* xics.vhdl:295:9  */
  assign n5390_o = n5387_o & n5389_o;
  /* xics.vhdl:295:9  */
  assign n5391_o = n5387_o & n5388_o;
  /* xics.vhdl:295:9  */
  assign n5392_o = n5386_o & n5389_o;
  /* xics.vhdl:295:9  */
  assign n5393_o = n5386_o & n5388_o;
  /* xics.vhdl:295:9  */
  assign n5394_o = n3408_o[0];
  /* xics.vhdl:295:9  */
  assign n5395_o = ~n5394_o;
  /* xics.vhdl:295:9  */
  assign n5396_o = n5390_o & n5395_o;
  /* xics.vhdl:295:9  */
  assign n5397_o = n5390_o & n5394_o;
  /* xics.vhdl:295:9  */
  assign n5398_o = n5391_o & n5395_o;
  /* xics.vhdl:295:9  */
  assign n5399_o = n5391_o & n5394_o;
  /* xics.vhdl:295:9  */
  assign n5400_o = n5392_o & n5395_o;
  /* xics.vhdl:295:9  */
  assign n5401_o = n5392_o & n5394_o;
  /* xics.vhdl:295:9  */
  assign n5402_o = n5393_o & n5395_o;
  /* xics.vhdl:295:9  */
  assign n5403_o = n5393_o & n5394_o;
  assign n5404_o = n3416_o[0];
  /* xics.vhdl:295:9  */
  assign n5405_o = n5396_o ? 1'b1 : n5404_o;
  assign n5406_o = n3416_o[1];
  /* xics.vhdl:295:9  */
  assign n5407_o = n5397_o ? 1'b1 : n5406_o;
  assign n5408_o = n3416_o[2];
  /* xics.vhdl:295:9  */
  assign n5409_o = n5398_o ? 1'b1 : n5408_o;
  assign n5410_o = n3416_o[3];
  /* xics.vhdl:295:9  */
  assign n5411_o = n5399_o ? 1'b1 : n5410_o;
  assign n5412_o = n3416_o[4];
  /* xics.vhdl:295:9  */
  assign n5413_o = n5400_o ? 1'b1 : n5412_o;
  assign n5414_o = n3416_o[5];
  /* xics.vhdl:295:9  */
  assign n5415_o = n5401_o ? 1'b1 : n5414_o;
  assign n5416_o = n3416_o[6];
  /* xics.vhdl:295:9  */
  assign n5417_o = n5402_o ? 1'b1 : n5416_o;
  assign n5418_o = n3416_o[7];
  /* xics.vhdl:295:9  */
  assign n5419_o = n5403_o ? 1'b1 : n5418_o;
  assign n5420_o = {n5419_o, n5417_o, n5415_o, n5413_o, n5411_o, n5409_o, n5407_o, n5405_o};
  /* xics.vhdl:295:9  */
  assign n5421_o = n3425_o[2];
  /* xics.vhdl:295:9  */
  assign n5422_o = ~n5421_o;
  /* xics.vhdl:295:9  */
  assign n5423_o = n3425_o[1];
  /* xics.vhdl:295:9  */
  assign n5424_o = ~n5423_o;
  /* xics.vhdl:295:9  */
  assign n5425_o = n5422_o & n5424_o;
  /* xics.vhdl:295:9  */
  assign n5426_o = n5422_o & n5423_o;
  /* xics.vhdl:295:9  */
  assign n5427_o = n5421_o & n5424_o;
  /* xics.vhdl:295:9  */
  assign n5428_o = n5421_o & n5423_o;
  /* xics.vhdl:295:9  */
  assign n5429_o = n3425_o[0];
  /* xics.vhdl:295:9  */
  assign n5430_o = ~n5429_o;
  /* xics.vhdl:295:9  */
  assign n5431_o = n5425_o & n5430_o;
  /* xics.vhdl:295:9  */
  assign n5432_o = n5425_o & n5429_o;
  /* xics.vhdl:295:9  */
  assign n5433_o = n5426_o & n5430_o;
  /* xics.vhdl:295:9  */
  assign n5434_o = n5426_o & n5429_o;
  /* xics.vhdl:295:9  */
  assign n5435_o = n5427_o & n5430_o;
  /* xics.vhdl:295:9  */
  assign n5436_o = n5427_o & n5429_o;
  /* xics.vhdl:295:9  */
  assign n5437_o = n5428_o & n5430_o;
  /* xics.vhdl:295:9  */
  assign n5438_o = n5428_o & n5429_o;
  assign n5439_o = n3433_o[0];
  /* xics.vhdl:295:9  */
  assign n5440_o = n5431_o ? 1'b1 : n5439_o;
  assign n5441_o = n3433_o[1];
  /* xics.vhdl:295:9  */
  assign n5442_o = n5432_o ? 1'b1 : n5441_o;
  assign n5443_o = n3433_o[2];
  /* xics.vhdl:295:9  */
  assign n5444_o = n5433_o ? 1'b1 : n5443_o;
  assign n5445_o = n3433_o[3];
  /* xics.vhdl:295:9  */
  assign n5446_o = n5434_o ? 1'b1 : n5445_o;
  assign n5447_o = n3433_o[4];
  /* xics.vhdl:295:9  */
  assign n5448_o = n5435_o ? 1'b1 : n5447_o;
  assign n5449_o = n3433_o[5];
  /* xics.vhdl:295:9  */
  assign n5450_o = n5436_o ? 1'b1 : n5449_o;
  assign n5451_o = n3433_o[6];
  /* xics.vhdl:295:9  */
  assign n5452_o = n5437_o ? 1'b1 : n5451_o;
  assign n5453_o = n3433_o[7];
  /* xics.vhdl:295:9  */
  assign n5454_o = n5438_o ? 1'b1 : n5453_o;
  assign n5455_o = {n5454_o, n5452_o, n5450_o, n5448_o, n5446_o, n5444_o, n5442_o, n5440_o};
  /* xics.vhdl:295:9  */
  assign n5456_o = n3442_o[2];
  /* xics.vhdl:295:9  */
  assign n5457_o = ~n5456_o;
  /* xics.vhdl:295:9  */
  assign n5458_o = n3442_o[1];
  /* xics.vhdl:295:9  */
  assign n5459_o = ~n5458_o;
  /* xics.vhdl:295:9  */
  assign n5460_o = n5457_o & n5459_o;
  /* xics.vhdl:295:9  */
  assign n5461_o = n5457_o & n5458_o;
  /* xics.vhdl:295:9  */
  assign n5462_o = n5456_o & n5459_o;
  /* xics.vhdl:295:9  */
  assign n5463_o = n5456_o & n5458_o;
  /* xics.vhdl:295:9  */
  assign n5464_o = n3442_o[0];
  /* xics.vhdl:295:9  */
  assign n5465_o = ~n5464_o;
  /* xics.vhdl:295:9  */
  assign n5466_o = n5460_o & n5465_o;
  /* xics.vhdl:295:9  */
  assign n5467_o = n5460_o & n5464_o;
  /* xics.vhdl:295:9  */
  assign n5468_o = n5461_o & n5465_o;
  /* xics.vhdl:295:9  */
  assign n5469_o = n5461_o & n5464_o;
  /* xics.vhdl:295:9  */
  assign n5470_o = n5462_o & n5465_o;
  /* xics.vhdl:295:9  */
  assign n5471_o = n5462_o & n5464_o;
  /* xics.vhdl:295:9  */
  assign n5472_o = n5463_o & n5465_o;
  /* xics.vhdl:295:9  */
  assign n5473_o = n5463_o & n5464_o;
  assign n5474_o = n3450_o[0];
  /* xics.vhdl:295:9  */
  assign n5475_o = n5466_o ? 1'b1 : n5474_o;
  assign n5476_o = n3450_o[1];
  /* xics.vhdl:295:9  */
  assign n5477_o = n5467_o ? 1'b1 : n5476_o;
  assign n5478_o = n3450_o[2];
  /* xics.vhdl:295:9  */
  assign n5479_o = n5468_o ? 1'b1 : n5478_o;
  assign n5480_o = n3450_o[3];
  /* xics.vhdl:295:9  */
  assign n5481_o = n5469_o ? 1'b1 : n5480_o;
  assign n5482_o = n3450_o[4];
  /* xics.vhdl:295:9  */
  assign n5483_o = n5470_o ? 1'b1 : n5482_o;
  assign n5484_o = n3450_o[5];
  /* xics.vhdl:295:9  */
  assign n5485_o = n5471_o ? 1'b1 : n5484_o;
  assign n5486_o = n3450_o[6];
  /* xics.vhdl:295:9  */
  assign n5487_o = n5472_o ? 1'b1 : n5486_o;
  assign n5488_o = n3450_o[7];
  /* xics.vhdl:295:9  */
  assign n5489_o = n5473_o ? 1'b1 : n5488_o;
  assign n5490_o = {n5489_o, n5487_o, n5485_o, n5483_o, n5481_o, n5479_o, n5477_o, n5475_o};
  /* xics.vhdl:295:9  */
  assign n5491_o = n3459_o[2];
  /* xics.vhdl:295:9  */
  assign n5492_o = ~n5491_o;
  /* xics.vhdl:295:9  */
  assign n5493_o = n3459_o[1];
  /* xics.vhdl:295:9  */
  assign n5494_o = ~n5493_o;
  /* xics.vhdl:295:9  */
  assign n5495_o = n5492_o & n5494_o;
  /* xics.vhdl:295:9  */
  assign n5496_o = n5492_o & n5493_o;
  /* xics.vhdl:295:9  */
  assign n5497_o = n5491_o & n5494_o;
  /* xics.vhdl:295:9  */
  assign n5498_o = n5491_o & n5493_o;
  /* xics.vhdl:295:9  */
  assign n5499_o = n3459_o[0];
  /* xics.vhdl:295:9  */
  assign n5500_o = ~n5499_o;
  /* xics.vhdl:295:9  */
  assign n5501_o = n5495_o & n5500_o;
  /* xics.vhdl:295:9  */
  assign n5502_o = n5495_o & n5499_o;
  /* xics.vhdl:295:9  */
  assign n5503_o = n5496_o & n5500_o;
  /* xics.vhdl:295:9  */
  assign n5504_o = n5496_o & n5499_o;
  /* xics.vhdl:295:9  */
  assign n5505_o = n5497_o & n5500_o;
  /* xics.vhdl:295:9  */
  assign n5506_o = n5497_o & n5499_o;
  /* xics.vhdl:295:9  */
  assign n5507_o = n5498_o & n5500_o;
  /* xics.vhdl:295:9  */
  assign n5508_o = n5498_o & n5499_o;
  assign n5509_o = n3467_o[0];
  /* xics.vhdl:295:9  */
  assign n5510_o = n5501_o ? 1'b1 : n5509_o;
  assign n5511_o = n3467_o[1];
  /* xics.vhdl:295:9  */
  assign n5512_o = n5502_o ? 1'b1 : n5511_o;
  assign n5513_o = n3467_o[2];
  /* xics.vhdl:295:9  */
  assign n5514_o = n5503_o ? 1'b1 : n5513_o;
  assign n5515_o = n3467_o[3];
  /* xics.vhdl:295:9  */
  assign n5516_o = n5504_o ? 1'b1 : n5515_o;
  assign n5517_o = n3467_o[4];
  /* xics.vhdl:295:9  */
  assign n5518_o = n5505_o ? 1'b1 : n5517_o;
  assign n5519_o = n3467_o[5];
  /* xics.vhdl:295:9  */
  assign n5520_o = n5506_o ? 1'b1 : n5519_o;
  assign n5521_o = n3467_o[6];
  /* xics.vhdl:295:9  */
  assign n5522_o = n5507_o ? 1'b1 : n5521_o;
  assign n5523_o = n3467_o[7];
  /* xics.vhdl:295:9  */
  assign n5524_o = n5508_o ? 1'b1 : n5523_o;
  assign n5525_o = {n5524_o, n5522_o, n5520_o, n5518_o, n5516_o, n5514_o, n5512_o, n5510_o};
  /* xics.vhdl:295:9  */
  assign n5526_o = n3476_o[2];
  /* xics.vhdl:295:9  */
  assign n5527_o = ~n5526_o;
  /* xics.vhdl:295:9  */
  assign n5528_o = n3476_o[1];
  /* xics.vhdl:295:9  */
  assign n5529_o = ~n5528_o;
  /* xics.vhdl:295:9  */
  assign n5530_o = n5527_o & n5529_o;
  /* xics.vhdl:295:9  */
  assign n5531_o = n5527_o & n5528_o;
  /* xics.vhdl:295:9  */
  assign n5532_o = n5526_o & n5529_o;
  /* xics.vhdl:295:9  */
  assign n5533_o = n5526_o & n5528_o;
  /* xics.vhdl:295:9  */
  assign n5534_o = n3476_o[0];
  /* xics.vhdl:295:9  */
  assign n5535_o = ~n5534_o;
  /* xics.vhdl:295:9  */
  assign n5536_o = n5530_o & n5535_o;
  /* xics.vhdl:295:9  */
  assign n5537_o = n5530_o & n5534_o;
  /* xics.vhdl:295:9  */
  assign n5538_o = n5531_o & n5535_o;
  /* xics.vhdl:295:9  */
  assign n5539_o = n5531_o & n5534_o;
  /* xics.vhdl:295:9  */
  assign n5540_o = n5532_o & n5535_o;
  /* xics.vhdl:295:9  */
  assign n5541_o = n5532_o & n5534_o;
  /* xics.vhdl:295:9  */
  assign n5542_o = n5533_o & n5535_o;
  /* xics.vhdl:295:9  */
  assign n5543_o = n5533_o & n5534_o;
  assign n5544_o = n3484_o[0];
  /* xics.vhdl:295:9  */
  assign n5545_o = n5536_o ? 1'b1 : n5544_o;
  assign n5546_o = n3484_o[1];
  /* xics.vhdl:295:9  */
  assign n5547_o = n5537_o ? 1'b1 : n5546_o;
  assign n5548_o = n3484_o[2];
  /* xics.vhdl:295:9  */
  assign n5549_o = n5538_o ? 1'b1 : n5548_o;
  assign n5550_o = n3484_o[3];
  /* xics.vhdl:295:9  */
  assign n5551_o = n5539_o ? 1'b1 : n5550_o;
  assign n5552_o = n3484_o[4];
  /* xics.vhdl:295:9  */
  assign n5553_o = n5540_o ? 1'b1 : n5552_o;
  assign n5554_o = n3484_o[5];
  /* xics.vhdl:295:9  */
  assign n5555_o = n5541_o ? 1'b1 : n5554_o;
  assign n5556_o = n3484_o[6];
  /* xics.vhdl:295:9  */
  assign n5557_o = n5542_o ? 1'b1 : n5556_o;
  assign n5558_o = n3484_o[7];
  /* xics.vhdl:295:9  */
  assign n5559_o = n5543_o ? 1'b1 : n5558_o;
  assign n5560_o = {n5559_o, n5557_o, n5555_o, n5553_o, n5551_o, n5549_o, n5547_o, n5545_o};
  /* xics.vhdl:295:9  */
  assign n5561_o = n3493_o[2];
  /* xics.vhdl:295:9  */
  assign n5562_o = ~n5561_o;
  /* xics.vhdl:295:9  */
  assign n5563_o = n3493_o[1];
  /* xics.vhdl:295:9  */
  assign n5564_o = ~n5563_o;
  /* xics.vhdl:295:9  */
  assign n5565_o = n5562_o & n5564_o;
  /* xics.vhdl:295:9  */
  assign n5566_o = n5562_o & n5563_o;
  /* xics.vhdl:295:9  */
  assign n5567_o = n5561_o & n5564_o;
  /* xics.vhdl:295:9  */
  assign n5568_o = n5561_o & n5563_o;
  /* xics.vhdl:295:9  */
  assign n5569_o = n3493_o[0];
  /* xics.vhdl:295:9  */
  assign n5570_o = ~n5569_o;
  /* xics.vhdl:295:9  */
  assign n5571_o = n5565_o & n5570_o;
  /* xics.vhdl:295:9  */
  assign n5572_o = n5565_o & n5569_o;
  /* xics.vhdl:295:9  */
  assign n5573_o = n5566_o & n5570_o;
  /* xics.vhdl:295:9  */
  assign n5574_o = n5566_o & n5569_o;
  /* xics.vhdl:295:9  */
  assign n5575_o = n5567_o & n5570_o;
  /* xics.vhdl:295:9  */
  assign n5576_o = n5567_o & n5569_o;
  /* xics.vhdl:295:9  */
  assign n5577_o = n5568_o & n5570_o;
  /* xics.vhdl:295:9  */
  assign n5578_o = n5568_o & n5569_o;
  assign n5579_o = n3501_o[0];
  /* xics.vhdl:295:9  */
  assign n5580_o = n5571_o ? 1'b1 : n5579_o;
  assign n5581_o = n3501_o[1];
  /* xics.vhdl:295:9  */
  assign n5582_o = n5572_o ? 1'b1 : n5581_o;
  assign n5583_o = n3501_o[2];
  /* xics.vhdl:295:9  */
  assign n5584_o = n5573_o ? 1'b1 : n5583_o;
  assign n5585_o = n3501_o[3];
  /* xics.vhdl:295:9  */
  assign n5586_o = n5574_o ? 1'b1 : n5585_o;
  assign n5587_o = n3501_o[4];
  /* xics.vhdl:295:9  */
  assign n5588_o = n5575_o ? 1'b1 : n5587_o;
  assign n5589_o = n3501_o[5];
  /* xics.vhdl:295:9  */
  assign n5590_o = n5576_o ? 1'b1 : n5589_o;
  assign n5591_o = n3501_o[6];
  /* xics.vhdl:295:9  */
  assign n5592_o = n5577_o ? 1'b1 : n5591_o;
  assign n5593_o = n3501_o[7];
  /* xics.vhdl:295:9  */
  assign n5594_o = n5578_o ? 1'b1 : n5593_o;
  assign n5595_o = {n5594_o, n5592_o, n5590_o, n5588_o, n5586_o, n5584_o, n5582_o, n5580_o};
  /* xics.vhdl:295:9  */
  assign n5596_o = n3510_o[2];
  /* xics.vhdl:295:9  */
  assign n5597_o = ~n5596_o;
  /* xics.vhdl:295:9  */
  assign n5598_o = n3510_o[1];
  /* xics.vhdl:295:9  */
  assign n5599_o = ~n5598_o;
  /* xics.vhdl:295:9  */
  assign n5600_o = n5597_o & n5599_o;
  /* xics.vhdl:295:9  */
  assign n5601_o = n5597_o & n5598_o;
  /* xics.vhdl:295:9  */
  assign n5602_o = n5596_o & n5599_o;
  /* xics.vhdl:295:9  */
  assign n5603_o = n5596_o & n5598_o;
  /* xics.vhdl:295:9  */
  assign n5604_o = n3510_o[0];
  /* xics.vhdl:295:9  */
  assign n5605_o = ~n5604_o;
  /* xics.vhdl:295:9  */
  assign n5606_o = n5600_o & n5605_o;
  /* xics.vhdl:295:9  */
  assign n5607_o = n5600_o & n5604_o;
  /* xics.vhdl:295:9  */
  assign n5608_o = n5601_o & n5605_o;
  /* xics.vhdl:295:9  */
  assign n5609_o = n5601_o & n5604_o;
  /* xics.vhdl:295:9  */
  assign n5610_o = n5602_o & n5605_o;
  /* xics.vhdl:295:9  */
  assign n5611_o = n5602_o & n5604_o;
  /* xics.vhdl:295:9  */
  assign n5612_o = n5603_o & n5605_o;
  /* xics.vhdl:295:9  */
  assign n5613_o = n5603_o & n5604_o;
  assign n5614_o = n3518_o[0];
  /* xics.vhdl:295:9  */
  assign n5615_o = n5606_o ? 1'b1 : n5614_o;
  assign n5616_o = n3518_o[1];
  /* xics.vhdl:295:9  */
  assign n5617_o = n5607_o ? 1'b1 : n5616_o;
  assign n5618_o = n3518_o[2];
  /* xics.vhdl:295:9  */
  assign n5619_o = n5608_o ? 1'b1 : n5618_o;
  assign n5620_o = n3518_o[3];
  /* xics.vhdl:295:9  */
  assign n5621_o = n5609_o ? 1'b1 : n5620_o;
  assign n5622_o = n3518_o[4];
  /* xics.vhdl:295:9  */
  assign n5623_o = n5610_o ? 1'b1 : n5622_o;
  assign n5624_o = n3518_o[5];
  /* xics.vhdl:295:9  */
  assign n5625_o = n5611_o ? 1'b1 : n5624_o;
  assign n5626_o = n3518_o[6];
  /* xics.vhdl:295:9  */
  assign n5627_o = n5612_o ? 1'b1 : n5626_o;
  assign n5628_o = n3518_o[7];
  /* xics.vhdl:295:9  */
  assign n5629_o = n5613_o ? 1'b1 : n5628_o;
  assign n5630_o = {n5629_o, n5627_o, n5625_o, n5623_o, n5621_o, n5619_o, n5617_o, n5615_o};
endmodule

module xics_icp
  (input  clk,
   input  rst,
   input  [29:0] wb_in_adr,
   input  [31:0] wb_in_dat,
   input  [3:0] wb_in_sel,
   input  wb_in_cyc,
   input  wb_in_stb,
   input  wb_in_we,
   input  [3:0] ics_in_src,
   input  [7:0] ics_in_pri,
   output [31:0] wb_out_dat,
   output wb_out_ack,
   output wb_out_stall,
   output core_irq_out);
  wire [68:0] n2897_o;
  wire [31:0] n2899_o;
  wire n2900_o;
  wire n2901_o;
  wire [11:0] n2902_o;
  wire [73:0] r;
  wire [73:0] r_next;
  wire n2906_o;
  wire [31:0] n2910_o;
  wire n2911_o;
  wire [31:0] n2922_o;
  wire [7:0] n2928_o;
  wire [7:0] n2931_o;
  wire [7:0] n2933_o;
  wire [7:0] n2935_o;
  wire [31:0] n2936_o;
  wire n2937_o;
  wire n2938_o;
  wire n2939_o;
  wire n2941_o;
  wire [5:0] n2942_o;
  wire [7:0] n2944_o;
  wire [7:0] n2945_o;
  wire n2947_o;
  wire [7:0] n2948_o;
  wire n2956_o;
  wire [7:0] n2957_o;
  wire n2965_o;
  wire [2:0] n2966_o;
  wire [7:0] n2967_o;
  reg [7:0] n2968_o;
  wire [7:0] n2969_o;
  reg [7:0] n2970_o;
  wire [5:0] n2971_o;
  wire [7:0] n2973_o;
  wire [7:0] n2974_o;
  wire [23:0] n2975_o;
  wire [31:0] n2976_o;
  wire n2978_o;
  wire [7:0] n2979_o;
  wire [23:0] n2980_o;
  wire [31:0] n2981_o;
  wire [3:0] n2982_o;
  wire n2984_o;
  wire n2987_o;
  wire n2989_o;
  wire [7:0] n2990_o;
  wire n2992_o;
  wire [2:0] n2993_o;
  reg n2995_o;
  wire [23:0] n2996_o;
  wire [23:0] n2997_o;
  reg [23:0] n2999_o;
  wire [7:0] n3000_o;
  wire [7:0] n3001_o;
  reg [7:0] n3003_o;
  wire [15:0] n3004_o;
  wire n3008_o;
  wire [31:0] n3009_o;
  wire [31:0] n3011_o;
  wire n3013_o;
  wire n3014_o;
  wire n3018_o;
  wire [31:0] n3021_o;
  wire [7:0] n3026_o;
  wire n3028_o;
  wire [3:0] n3029_o;
  wire [23:0] n3031_o;
  wire [7:0] n3032_o;
  wire [23:0] n3033_o;
  wire [7:0] n3035_o;
  wire [7:0] n3037_o;
  wire n3038_o;
  wire [7:0] n3040_o;
  wire [23:0] n3041_o;
  wire [7:0] n3042_o;
  wire [7:0] n3043_o;
  wire [7:0] n3044_o;
  wire [7:0] n3045_o;
  wire [7:0] n3046_o;
  wire [7:0] n3047_o;
  wire [7:0] n3048_o;
  wire [7:0] n3049_o;
  wire [7:0] n3056_o;
  wire [7:0] n3059_o;
  wire [7:0] n3061_o;
  wire [7:0] n3063_o;
  wire [31:0] n3064_o;
  wire [73:0] n3065_o;
  wire [7:0] n3066_o;
  wire n3067_o;
  wire n3072_o;
  wire [73:0] n3074_o;
  wire [73:0] n3075_o;
  reg [73:0] n3078_q;
  wire [33:0] n3079_o;
  reg n3080_q;
  assign wb_out_dat = n2899_o;
  assign wb_out_ack = n2900_o;
  assign wb_out_stall = n2901_o;
  assign core_irq_out = n3080_q;
  /* spi_flash_ctrl.vhdl:154:23  */
  assign n2897_o = {wb_in_we, wb_in_stb, wb_in_cyc, wb_in_sel, wb_in_dat, wb_in_adr};
  /* spi_flash_ctrl.vhdl:152:27  */
  assign n2899_o = n3079_o[31:0];
  /* spi_flash_ctrl.vhdl:151:24  */
  assign n2900_o = n3079_o[32];
  /* spi_flash_ctrl.vhdl:150:24  */
  assign n2901_o = n3079_o[33];
  /* spi_flash_ctrl.vhdl:146:28  */
  assign n2902_o = {ics_in_pri, ics_in_src};
  /* xics.vhdl:55:12  */
  assign r = n3078_q; // (signal)
  /* xics.vhdl:55:15  */
  assign r_next = n3075_o; // (signal)
  /* xics.vhdl:71:31  */
  assign n2906_o = r[40];
  /* xics.vhdl:75:21  */
  assign n2910_o = r[72:41];
  /* xics.vhdl:76:21  */
  assign n2911_o = r[73];
  /* xics.vhdl:104:30  */
  assign n2922_o = n2897_o[61:30];
  /* xics.vhdl:86:33  */
  assign n2928_o = n2922_o[31:24];
  /* xics.vhdl:87:33  */
  assign n2931_o = n2922_o[23:16];
  /* xics.vhdl:88:33  */
  assign n2933_o = n2922_o[15:8];
  /* xics.vhdl:89:33  */
  assign n2935_o = n2922_o[7:0];
  /* spi_flash_ctrl.vhdl:574:18  */
  assign n2936_o = {n2935_o, n2933_o, n2931_o, n2928_o};
  /* xics.vhdl:107:18  */
  assign n2937_o = n2897_o[66];
  /* xics.vhdl:107:38  */
  assign n2938_o = n2897_o[67];
  /* xics.vhdl:107:28  */
  assign n2939_o = n2937_o & n2938_o;
  /* xics.vhdl:109:22  */
  assign n2941_o = n2897_o[68];
  /* xics.vhdl:111:31  */
  assign n2942_o = n2897_o[5:0];
  /* xics.vhdl:111:44  */
  assign n2944_o = {n2942_o, 2'b00};
  /* xics.vhdl:114:36  */
  assign n2945_o = n2936_o[31:24];
  /* xics.vhdl:112:17  */
  assign n2947_o = n2944_o == 8'b00000000;
  /* xics.vhdl:116:36  */
  assign n2948_o = n2936_o[31:24];
  /* xics.vhdl:115:17  */
  assign n2956_o = n2944_o == 8'b00000100;
  /* xics.vhdl:125:36  */
  assign n2957_o = n2936_o[31:24];
  /* xics.vhdl:124:17  */
  assign n2965_o = n2944_o == 8'b00001100;
  assign n2966_o = {n2965_o, n2956_o, n2947_o};
  assign n2967_o = r[31:24];
  /* xics.vhdl:111:17  */
  always @*
    case (n2966_o)
      3'b100: n2968_o = n2967_o;
      3'b010: n2968_o = n2948_o;
      3'b001: n2968_o = n2945_o;
      default: n2968_o = n2967_o;
    endcase
  assign n2969_o = r[39:32];
  /* xics.vhdl:111:17  */
  always @*
    case (n2966_o)
      3'b100: n2970_o = n2957_o;
      3'b010: n2970_o = n2969_o;
      3'b001: n2970_o = n2969_o;
      default: n2970_o = n2969_o;
    endcase
  /* xics.vhdl:138:31  */
  assign n2971_o = n2897_o[5:0];
  /* xics.vhdl:138:44  */
  assign n2973_o = {n2971_o, 2'b00};
  /* xics.vhdl:141:33  */
  assign n2974_o = r[31:24];
  /* xics.vhdl:141:42  */
  assign n2975_o = r[23:0];
  /* xics.vhdl:141:38  */
  assign n2976_o = {n2974_o, n2975_o};
  /* xics.vhdl:139:17  */
  assign n2978_o = n2973_o == 8'b00000000;
  /* xics.vhdl:144:33  */
  assign n2979_o = r[31:24];
  /* xics.vhdl:144:42  */
  assign n2980_o = r[23:0];
  /* xics.vhdl:144:38  */
  assign n2981_o = {n2979_o, n2980_o};
  /* xics.vhdl:145:30  */
  assign n2982_o = n2897_o[65:62];
  /* xics.vhdl:145:34  */
  assign n2984_o = n2982_o == 4'b1111;
  /* xics.vhdl:145:21  */
  assign n2987_o = n2984_o ? 1'b1 : 1'b0;
  /* xics.vhdl:142:17  */
  assign n2989_o = n2973_o == 8'b00000100;
  /* xics.vhdl:150:47  */
  assign n2990_o = r[39:32];
  /* xics.vhdl:148:17  */
  assign n2992_o = n2973_o == 8'b00001100;
  assign n2993_o = {n2992_o, n2989_o, n2978_o};
  /* xics.vhdl:138:17  */
  always @*
    case (n2993_o)
      3'b100: n2995_o = 1'b0;
      3'b010: n2995_o = n2987_o;
      3'b001: n2995_o = 1'b0;
      default: n2995_o = 1'b0;
    endcase
  /* spi_flash_ctrl.vhdl:281:9  */
  assign n2996_o = n2976_o[23:0];
  /* spi_flash_ctrl.vhdl:273:5  */
  assign n2997_o = n2981_o[23:0];
  /* xics.vhdl:138:17  */
  always @*
    case (n2993_o)
      3'b100: n2999_o = 24'b000000000000000000000000;
      3'b010: n2999_o = n2997_o;
      3'b001: n2999_o = n2996_o;
      default: n2999_o = 24'b000000000000000000000000;
    endcase
  assign n3000_o = n2976_o[31:24];
  /* spi_flash_ctrl.vhdl:217:28  */
  assign n3001_o = n2981_o[31:24];
  /* xics.vhdl:138:17  */
  always @*
    case (n2993_o)
      3'b100: n3003_o = n2990_o;
      3'b010: n3003_o = n3001_o;
      3'b001: n3003_o = n3000_o;
      default: n3003_o = 8'b00000000;
    endcase
  assign n3004_o = {n2970_o, n2968_o};
  /* xics.vhdl:109:13  */
  assign n3008_o = n2941_o ? 1'b0 : n2995_o;
  assign n3009_o = {n3003_o, n2999_o};
  /* xics.vhdl:109:13  */
  assign n3011_o = n2941_o ? 32'b00000000000000000000000000000000 : n3009_o;
  /* xics.vhdl:107:9  */
  assign n3013_o = n2939_o & n2941_o;
  /* xics.vhdl:107:9  */
  assign n3014_o = n2939_o ? 1'b1 : 1'b0;
  /* xics.vhdl:107:9  */
  assign n3018_o = n2939_o ? n3008_o : 1'b0;
  /* xics.vhdl:107:9  */
  assign n3021_o = n2939_o ? n3011_o : 32'b00000000000000000000000000000000;
  /* xics.vhdl:160:19  */
  assign n3026_o = n2902_o[11:4];
  /* xics.vhdl:160:23  */
  assign n3028_o = n3026_o != 8'b11111111;
  /* xics.vhdl:161:41  */
  assign n3029_o = n2902_o[3:0];
  /* xics.vhdl:161:32  */
  assign n3031_o = {20'b00000000000000000001, n3029_o};
  /* xics.vhdl:162:40  */
  assign n3032_o = n2902_o[11:4];
  /* xics.vhdl:160:9  */
  assign n3033_o = n3028_o ? n3031_o : 24'b000000000000000000000000;
  /* xics.vhdl:160:9  */
  assign n3035_o = n3028_o ? n3032_o : 8'b11111111;
  /* xics.vhdl:166:23  */
  assign n3037_o = r[39:32];
  /* xics.vhdl:166:29  */
  assign n3038_o = $unsigned(n3037_o) < $unsigned(n3035_o);
  /* xics.vhdl:168:35  */
  assign n3040_o = r[39:32];
  /* xics.vhdl:166:9  */
  assign n3041_o = n3038_o ? 24'b000000000000000000000010 : n3033_o;
  /* xics.vhdl:166:9  */
  assign n3042_o = n3038_o ? n3040_o : n3035_o;
  assign n3043_o = n3004_o[7:0];
  assign n3044_o = r[31:24];
  /* xics.vhdl:107:9  */
  assign n3045_o = n3013_o ? n3043_o : n3044_o;
  /* xics.vhdl:172:9  */
  assign n3046_o = n3018_o ? n3042_o : n3045_o;
  assign n3047_o = n3004_o[15:8];
  assign n3048_o = r[39:32];
  /* xics.vhdl:107:9  */
  assign n3049_o = n3013_o ? n3047_o : n3048_o;
  /* xics.vhdl:86:33  */
  assign n3056_o = n3021_o[31:24];
  /* xics.vhdl:87:33  */
  assign n3059_o = n3021_o[23:16];
  /* xics.vhdl:88:33  */
  assign n3061_o = n3021_o[15:8];
  /* xics.vhdl:89:33  */
  assign n3063_o = n3021_o[7:0];
  assign n3064_o = {n3063_o, n3061_o, n3059_o, n3056_o};
  assign n3065_o = {n3014_o, n3064_o, 1'b0, n3049_o, n3046_o, n3041_o};
  /* xics.vhdl:182:52  */
  assign n3066_o = n3065_o[31:24];
  /* xics.vhdl:182:39  */
  assign n3067_o = $unsigned(n3042_o) < $unsigned(n3066_o);
  /* xics.vhdl:182:9  */
  assign n3072_o = n3067_o ? 1'b1 : 1'b0;
  assign n3074_o = {n3014_o, n3064_o, n3072_o, n3049_o, n3046_o, n3041_o};
  /* xics.vhdl:191:9  */
  assign n3075_o = rst ? 74'b00000000000000000000000000000000001111111100000000000000000000000000000000 : n3074_o;
  /* xics.vhdl:67:9  */
  always @(posedge clk)
    n3078_q <= r_next;
  /* xics.vhdl:67:9  */
  assign n3079_o = {1'b0, n2911_o, n2910_o};
  /* xics.vhdl:67:9  */
  always @(posedge clk)
    n3080_q <= n2906_o;
endmodule

module spi_flash_ctrl_4_4_1489f923c4dca729178b3e3233458550d8dddf29
  (input  clk,
   input  rst,
   input  [29:0] wb_in_adr,
   input  [31:0] wb_in_dat,
   input  [3:0] wb_in_sel,
   input  wb_in_cyc,
   input  wb_in_stb,
   input  wb_in_we,
   input  wb_sel_reg,
   input  wb_sel_map,
   input  [3:0] sdat_i,
   output [31:0] wb_out_dat,
   output wb_out_ack,
   output wb_out_stall,
   output sck,
   output cs_n,
   output [3:0] sdat_o,
   output [3:0] sdat_oe);
  wire [68:0] n2023_o;
  wire [31:0] n2025_o;
  wire n2026_o;
  wire n2027_o;
  reg [15:0] ctrl_reg;
  reg [29:0] auto_cfg_reg;
  wire cmd_valid;
  wire [7:0] cmd_clk_div;
  wire [2:0] cmd_mode;
  wire cmd_ready;
  wire [2:0] d_clks;
  wire [7:0] d_rx;
  wire [7:0] d_tx;
  wire d_ack;
  wire bus_idle;
  wire pending_read;
  wire [68:0] wb_req;
  wire [68:0] wb_stash;
  wire [33:0] wb_rsp;
  wire wb_valid;
  wire wb_reg_valid;
  wire wb_reg_dat_v;
  wire wb_map_valid;
  wire [2:0] wb_reg;
  wire auto_cs;
  wire auto_cmd_valid;
  wire [2:0] auto_cmd_mode;
  wire [7:0] auto_d_txd;
  wire [2:0] auto_d_clks;
  wire [31:0] auto_data_next;
  wire [5:0] auto_cnt_next;
  wire auto_ack;
  wire [4:0] auto_next;
  wire [31:0] auto_lad_next;
  wire auto_latch_adr;
  reg [31:0] auto_data;
  reg [5:0] auto_cnt;
  reg [4:0] auto_state;
  wire [31:0] auto_last_addr;
  wire spi_rxtx_cmd_ready_o;
  wire [7:0] spi_rxtx_d_rxd_o;
  wire spi_rxtx_d_ack_o;
  wire spi_rxtx_bus_idle_o;
  wire spi_rxtx_sck;
  wire [3:0] spi_rxtx_sdat_o;
  wire [3:0] spi_rxtx_sdat_oe;
  wire n2044_o;
  wire n2045_o;
  wire n2046_o;
  wire n2047_o;
  wire n2048_o;
  wire [2:0] n2049_o;
  wire [2:0] n2050_o;
  wire n2054_o;
  wire n2055_o;
  wire n2059_o;
  wire n2060_o;
  wire n2061_o;
  wire n2063_o;
  wire n2064_o;
  wire n2068_o;
  wire n2069_o;
  wire n2070_o;
  wire n2071_o;
  wire n2072_o;
  wire [7:0] n2073_o;
  wire [3:0] n2075_o;
  wire n2077_o;
  wire n2078_o;
  wire [2:0] n2080_o;
  wire [3:0] n2081_o;
  wire n2083_o;
  wire n2084_o;
  wire [2:0] n2086_o;
  wire n2087_o;
  wire [2:0] n2089_o;
  wire [2:0] n2090_o;
  wire [2:0] n2093_o;
  wire [2:0] n2094_o;
  wire [2:0] n2096_o;
  wire [7:0] n2097_o;
  wire n2098_o;
  wire n2099_o;
  wire [7:0] n2100_o;
  wire n2102_o;
  wire n2103_o;
  wire n2104_o;
  wire [7:0] n2105_o;
  wire [2:0] n2106_o;
  wire [2:0] n2107_o;
  wire [7:0] n2108_o;
  wire n2118_o;
  wire n2119_o;
  wire n2120_o;
  wire n2121_o;
  wire n2122_o;
  wire n2123_o;
  wire n2124_o;
  wire n2125_o;
  wire n2127_o;
  wire n2128_o;
  wire [32:0] n2129_o;
  wire [68:0] n2130_o;
  wire n2131_o;
  wire n2132_o;
  wire n2133_o;
  wire n2135_o;
  wire n2136_o;
  wire n2137_o;
  wire [1:0] n2138_o;
  wire [65:0] n2139_o;
  wire [65:0] n2140_o;
  wire [65:0] n2141_o;
  wire [1:0] n2142_o;
  wire [1:0] n2143_o;
  wire n2144_o;
  wire n2145_o;
  wire n2146_o;
  wire n2147_o;
  wire [68:0] n2148_o;
  wire [68:0] n2149_o;
  wire n2150_o;
  wire [68:0] n2151_o;
  wire [33:0] n2152_o;
  wire [1:0] n2153_o;
  wire [31:0] n2154_o;
  wire [31:0] n2155_o;
  wire [31:0] n2156_o;
  wire [1:0] n2157_o;
  wire [1:0] n2158_o;
  wire [68:0] n2159_o;
  wire [6:0] n2160_o;
  wire [61:0] n2161_o;
  wire [61:0] n2162_o;
  wire [61:0] n2163_o;
  wire [6:0] n2164_o;
  wire [6:0] n2165_o;
  wire [33:0] n2166_o;
  wire [68:0] n2169_o;
  wire [15:0] n2175_o;
  wire [23:0] n2176_o;
  wire [31:0] n2177_o;
  wire n2179_o;
  wire n2180_o;
  wire n2182_o;
  wire n2183_o;
  wire n2184_o;
  wire n2185_o;
  wire n2187_o;
  wire n2188_o;
  wire n2189_o;
  wire [1:0] n2190_o;
  wire n2191_o;
  wire n2192_o;
  wire n2193_o;
  wire n2194_o;
  wire n2196_o;
  wire n2197_o;
  wire [3:0] n2216_o;
  wire [3:0] n2217_o;
  wire [3:0] n2218_o;
  wire [3:0] n2219_o;
  wire [15:0] n2220_o;
  wire [31:0] n2221_o;
  wire n2223_o;
  wire [31:0] n2226_o;
  wire n2228_o;
  wire [1:0] n2229_o;
  reg [31:0] n2230_o;
  wire [33:0] n2232_o;
  wire [32:0] n2233_o;
  wire [32:0] n2234_o;
  wire [32:0] n2235_o;
  wire n2236_o;
  wire n2237_o;
  wire [33:0] n2238_o;
  wire [33:0] n2239_o;
  wire [33:0] n2240_o;
  wire [1:0] n2241_o;
  wire [31:0] n2242_o;
  wire [31:0] n2243_o;
  wire [1:0] n2244_o;
  wire [1:0] n2245_o;
  wire [33:0] n2246_o;
  wire [33:0] n2247_o;
  wire n2249_o;
  wire n2250_o;
  wire n2252_o;
  wire n2253_o;
  wire n2254_o;
  wire n2255_o;
  wire n2256_o;
  wire n2257_o;
  wire n2258_o;
  wire [31:0] n2259_o;
  wire [31:0] n2260_o;
  wire [31:0] n2261_o;
  wire [31:0] n2265_o;
  wire [31:0] n2266_o;
  wire [5:0] n2267_o;
  wire [4:0] n2269_o;
  wire [31:0] n2271_o;
  wire [27:0] n2280_o;
  wire [29:0] n2282_o;
  wire [31:0] n2284_o;
  wire [31:0] n2286_o;
  wire n2287_o;
  wire n2288_o;
  wire n2289_o;
  wire [31:0] n2290_o;
  wire n2292_o;
  wire [31:0] n2293_o;
  wire [31:0] n2295_o;
  wire [5:0] n2296_o;
  wire [5:0] n2297_o;
  wire n2299_o;
  wire n2301_o;
  wire n2302_o;
  wire n2304_o;
  wire n2305_o;
  wire n2308_o;
  wire n2310_o;
  wire n2311_o;
  wire n2312_o;
  wire n2313_o;
  wire n2314_o;
  wire [5:0] n2316_o;
  wire n2319_o;
  wire [4:0] n2321_o;
  wire [5:0] n2322_o;
  wire n2324_o;
  wire [4:0] n2325_o;
  wire n2327_o;
  wire [31:0] n2328_o;
  wire n2330_o;
  wire [4:0] n2332_o;
  wire n2334_o;
  wire [7:0] n2335_o;
  wire n2336_o;
  wire [4:0] n2339_o;
  wire [4:0] n2340_o;
  wire n2342_o;
  wire [7:0] n2343_o;
  wire [4:0] n2345_o;
  wire n2347_o;
  wire [7:0] n2348_o;
  wire [4:0] n2350_o;
  wire n2352_o;
  wire [7:0] n2353_o;
  wire [4:0] n2355_o;
  wire n2357_o;
  wire [7:0] n2358_o;
  wire [2:0] n2360_o;
  wire n2361_o;
  wire [4:0] n2364_o;
  wire [4:0] n2365_o;
  wire n2367_o;
  wire [2:0] n2368_o;
  wire [4:0] n2370_o;
  wire n2372_o;
  wire [1:0] n2373_o;
  wire [2:0] n2375_o;
  wire [1:0] n2382_o;
  wire n2383_o;
  wire [1:0] n2386_o;
  wire n2387_o;
  wire [2:0] n2390_o;
  wire [2:0] n2391_o;
  wire [4:0] n2393_o;
  wire n2395_o;
  wire [7:0] n2396_o;
  wire [7:0] n2397_o;
  wire [4:0] n2399_o;
  wire n2401_o;
  wire [1:0] n2402_o;
  wire [2:0] n2404_o;
  wire [1:0] n2411_o;
  wire n2412_o;
  wire [1:0] n2415_o;
  wire n2416_o;
  wire [2:0] n2419_o;
  wire [2:0] n2420_o;
  wire [4:0] n2422_o;
  wire n2424_o;
  wire [7:0] n2425_o;
  wire [7:0] n2426_o;
  wire [4:0] n2428_o;
  wire n2430_o;
  wire [1:0] n2431_o;
  wire [2:0] n2433_o;
  wire [1:0] n2440_o;
  wire n2441_o;
  wire [1:0] n2444_o;
  wire n2445_o;
  wire [2:0] n2448_o;
  wire [2:0] n2449_o;
  wire [4:0] n2451_o;
  wire n2453_o;
  wire [7:0] n2454_o;
  wire [7:0] n2455_o;
  wire [4:0] n2457_o;
  wire n2459_o;
  wire [1:0] n2460_o;
  wire [2:0] n2462_o;
  wire [1:0] n2469_o;
  wire n2470_o;
  wire [1:0] n2473_o;
  wire n2474_o;
  wire [2:0] n2477_o;
  wire [2:0] n2478_o;
  wire [4:0] n2480_o;
  wire n2482_o;
  wire [7:0] n2483_o;
  wire [7:0] n2484_o;
  wire [4:0] n2486_o;
  wire n2489_o;
  wire n2491_o;
  wire [5:0] n2492_o;
  wire n2495_o;
  wire n2496_o;
  wire n2497_o;
  wire n2498_o;
  wire n2499_o;
  wire n2500_o;
  wire [31:0] n2501_o;
  wire n2503_o;
  wire n2504_o;
  wire [5:0] n2506_o;
  wire [4:0] n2508_o;
  wire [5:0] n2509_o;
  wire [4:0] n2511_o;
  wire n2513_o;
  wire [31:0] n2514_o;
  wire n2516_o;
  wire [4:0] n2518_o;
  wire n2520_o;
  wire [19:0] n2521_o;
  reg n2534_o;
  reg [2:0] n2537_o;
  reg [7:0] n2540_o;
  reg [2:0] n2543_o;
  wire [7:0] n2544_o;
  reg [7:0] n2546_o;
  wire [7:0] n2547_o;
  reg [7:0] n2549_o;
  wire [7:0] n2550_o;
  reg [7:0] n2552_o;
  wire [7:0] n2553_o;
  reg [7:0] n2555_o;
  reg [5:0] n2557_o;
  reg n2561_o;
  reg [4:0] n2565_o;
  reg n2568_o;
  wire n2570_o;
  wire n2573_o;
  wire [2:0] n2576_o;
  wire [7:0] n2579_o;
  wire [2:0] n2582_o;
  wire [31:0] n2584_o;
  wire [31:0] n2585_o;
  wire [5:0] n2587_o;
  wire n2589_o;
  wire [4:0] n2592_o;
  wire n2594_o;
  wire n2599_o;
  wire n2600_o;
  wire [3:0] n2614_o;
  wire [3:0] n2615_o;
  wire [3:0] n2616_o;
  wire [7:0] n2617_o;
  wire [7:0] n2618_o;
  wire [29:0] n2619_o;
  wire [29:0] n2620_o;
  wire n2621_o;
  wire n2622_o;
  wire n2624_o;
  wire n2625_o;
  wire n2626_o;
  wire n2628_o;
  wire n2637_o;
  wire n2638_o;
  wire n2639_o;
  wire n2640_o;
  wire n2642_o;
  wire n2643_o;
  wire n2644_o;
  wire n2645_o;
  wire n2647_o;
  wire n2648_o;
  wire n2649_o;
  wire n2650_o;
  wire n2652_o;
  wire n2653_o;
  wire n2654_o;
  wire n2655_o;
  wire n2657_o;
  wire n2658_o;
  wire n2659_o;
  wire n2660_o;
  wire n2662_o;
  wire n2663_o;
  wire n2664_o;
  wire n2665_o;
  wire n2667_o;
  wire n2668_o;
  wire n2669_o;
  wire n2670_o;
  wire n2672_o;
  wire n2673_o;
  wire n2674_o;
  wire n2675_o;
  wire n2677_o;
  wire n2678_o;
  wire n2679_o;
  wire n2680_o;
  wire n2682_o;
  wire n2683_o;
  wire n2684_o;
  wire n2685_o;
  wire n2687_o;
  wire n2688_o;
  wire n2689_o;
  wire n2690_o;
  wire n2692_o;
  wire n2693_o;
  wire n2694_o;
  wire n2695_o;
  wire n2697_o;
  wire n2698_o;
  wire n2699_o;
  wire n2700_o;
  wire n2702_o;
  wire n2703_o;
  wire n2704_o;
  wire n2705_o;
  wire n2707_o;
  wire n2708_o;
  wire n2709_o;
  wire n2710_o;
  wire n2711_o;
  wire n2712_o;
  wire n2713_o;
  wire n2714_o;
  wire [15:0] n2715_o;
  wire [3:0] n2716_o;
  wire [15:0] n2717_o;
  wire [15:0] n2718_o;
  wire n2720_o;
  wire n2729_o;
  wire n2730_o;
  wire n2731_o;
  wire n2732_o;
  wire n2734_o;
  wire n2735_o;
  wire n2736_o;
  wire n2737_o;
  wire n2739_o;
  wire n2740_o;
  wire n2741_o;
  wire n2742_o;
  wire n2744_o;
  wire n2745_o;
  wire n2746_o;
  wire n2747_o;
  wire n2749_o;
  wire n2750_o;
  wire n2751_o;
  wire n2752_o;
  wire n2754_o;
  wire n2755_o;
  wire n2756_o;
  wire n2757_o;
  wire n2759_o;
  wire n2760_o;
  wire n2761_o;
  wire n2762_o;
  wire n2764_o;
  wire n2765_o;
  wire n2766_o;
  wire n2767_o;
  wire n2769_o;
  wire n2770_o;
  wire n2771_o;
  wire n2772_o;
  wire n2774_o;
  wire n2775_o;
  wire n2776_o;
  wire n2777_o;
  wire n2779_o;
  wire n2780_o;
  wire n2781_o;
  wire n2782_o;
  wire n2784_o;
  wire n2785_o;
  wire n2786_o;
  wire n2787_o;
  wire n2789_o;
  wire n2790_o;
  wire n2791_o;
  wire n2792_o;
  wire n2794_o;
  wire n2795_o;
  wire n2796_o;
  wire n2797_o;
  wire n2799_o;
  wire n2800_o;
  wire n2801_o;
  wire n2802_o;
  wire n2804_o;
  wire n2805_o;
  wire n2806_o;
  wire n2807_o;
  wire n2809_o;
  wire n2810_o;
  wire n2811_o;
  wire n2812_o;
  wire n2814_o;
  wire n2815_o;
  wire n2816_o;
  wire n2817_o;
  wire n2819_o;
  wire n2820_o;
  wire n2821_o;
  wire n2822_o;
  wire n2824_o;
  wire n2825_o;
  wire n2826_o;
  wire n2827_o;
  wire n2829_o;
  wire n2830_o;
  wire n2831_o;
  wire n2832_o;
  wire n2834_o;
  wire n2835_o;
  wire n2836_o;
  wire n2837_o;
  wire n2839_o;
  wire n2840_o;
  wire n2841_o;
  wire n2842_o;
  wire n2844_o;
  wire n2845_o;
  wire n2846_o;
  wire n2847_o;
  wire n2849_o;
  wire n2850_o;
  wire n2851_o;
  wire n2852_o;
  wire n2854_o;
  wire n2855_o;
  wire n2856_o;
  wire n2857_o;
  wire n2859_o;
  wire n2860_o;
  wire n2861_o;
  wire n2862_o;
  wire n2864_o;
  wire n2865_o;
  wire n2866_o;
  wire n2867_o;
  wire n2869_o;
  wire n2870_o;
  wire n2871_o;
  wire n2872_o;
  wire n2873_o;
  wire n2874_o;
  wire n2875_o;
  wire n2876_o;
  wire [29:0] n2877_o;
  wire [29:0] n2878_o;
  wire [3:0] n2879_o;
  wire [15:0] n2880_o;
  wire [15:0] n2881_o;
  wire n2882_o;
  reg [15:0] n2886_q;
  reg [29:0] n2887_q;
  reg n2888_q;
  reg [68:0] n2889_q;
  reg [68:0] n2890_q;
  wire [33:0] n2891_o;
  reg [31:0] n2892_q;
  reg [5:0] n2893_q;
  reg [4:0] n2894_q;
  reg [31:0] n2895_q;
  reg [33:0] n2896_q;
  assign wb_out_dat = n2025_o;
  assign wb_out_ack = n2026_o;
  assign wb_out_stall = n2027_o;
  assign sck = spi_rxtx_sck;
  assign cs_n = n2103_o;
  assign sdat_o = spi_rxtx_sdat_o;
  assign sdat_oe = spi_rxtx_sdat_oe;
  /* syscon.vhdl:35:9  */
  assign n2023_o = {wb_in_we, wb_in_stb, wb_in_cyc, wb_in_sel, wb_in_dat, wb_in_adr};
  /* syscon.vhdl:31:9  */
  assign n2025_o = n2896_q[31:0];
  assign n2026_o = n2896_q[32];
  /* syscon.vhdl:206:17  */
  assign n2027_o = n2896_q[33];
  /* spi_flash_ctrl.vhdl:53:12  */
  always @*
    ctrl_reg = n2886_q; // (isignal)
  initial
    ctrl_reg = 16'b0000000000000000;
  /* spi_flash_ctrl.vhdl:61:12  */
  always @*
    auto_cfg_reg = n2887_q; // (isignal)
  initial
    auto_cfg_reg = 30'b000000000000000000000000000000;
  /* spi_flash_ctrl.vhdl:77:12  */
  assign cmd_valid = n2104_o; // (signal)
  /* spi_flash_ctrl.vhdl:78:12  */
  assign cmd_clk_div = n2105_o; // (signal)
  /* spi_flash_ctrl.vhdl:79:12  */
  assign cmd_mode = n2106_o; // (signal)
  /* spi_flash_ctrl.vhdl:80:12  */
  assign cmd_ready = spi_rxtx_cmd_ready_o; // (signal)
  /* spi_flash_ctrl.vhdl:81:12  */
  assign d_clks = n2107_o; // (signal)
  /* spi_flash_ctrl.vhdl:82:12  */
  assign d_rx = spi_rxtx_d_rxd_o; // (signal)
  /* spi_flash_ctrl.vhdl:83:12  */
  assign d_tx = n2108_o; // (signal)
  /* spi_flash_ctrl.vhdl:84:12  */
  assign d_ack = spi_rxtx_d_ack_o; // (signal)
  /* spi_flash_ctrl.vhdl:85:12  */
  assign bus_idle = spi_rxtx_bus_idle_o; // (signal)
  /* spi_flash_ctrl.vhdl:88:12  */
  assign pending_read = n2888_q; // (signal)
  /* spi_flash_ctrl.vhdl:91:12  */
  assign wb_req = n2889_q; // (signal)
  /* spi_flash_ctrl.vhdl:92:12  */
  assign wb_stash = n2890_q; // (signal)
  /* spi_flash_ctrl.vhdl:93:12  */
  assign wb_rsp = n2891_o; // (signal)
  /* spi_flash_ctrl.vhdl:96:12  */
  assign wb_valid = n2046_o; // (signal)
  /* spi_flash_ctrl.vhdl:97:12  */
  assign wb_reg_valid = n2047_o; // (signal)
  /* spi_flash_ctrl.vhdl:98:12  */
  assign wb_reg_dat_v = n2055_o; // (signal)
  /* spi_flash_ctrl.vhdl:99:12  */
  assign wb_map_valid = n2048_o; // (signal)
  /* spi_flash_ctrl.vhdl:100:12  */
  assign wb_reg = n2050_o; // (signal)
  /* spi_flash_ctrl.vhdl:116:12  */
  assign auto_cs = n2570_o; // (signal)
  /* spi_flash_ctrl.vhdl:117:12  */
  assign auto_cmd_valid = n2573_o; // (signal)
  /* spi_flash_ctrl.vhdl:118:12  */
  assign auto_cmd_mode = n2576_o; // (signal)
  /* spi_flash_ctrl.vhdl:119:12  */
  assign auto_d_txd = n2579_o; // (signal)
  /* spi_flash_ctrl.vhdl:120:12  */
  assign auto_d_clks = n2582_o; // (signal)
  /* spi_flash_ctrl.vhdl:121:12  */
  assign auto_data_next = n2585_o; // (signal)
  /* spi_flash_ctrl.vhdl:122:12  */
  assign auto_cnt_next = n2587_o; // (signal)
  /* spi_flash_ctrl.vhdl:123:12  */
  assign auto_ack = n2589_o; // (signal)
  /* spi_flash_ctrl.vhdl:124:12  */
  assign auto_next = n2592_o; // (signal)
  /* spi_flash_ctrl.vhdl:125:12  */
  assign auto_lad_next = n2286_o; // (signal)
  /* spi_flash_ctrl.vhdl:126:12  */
  assign auto_latch_adr = n2594_o; // (signal)
  /* spi_flash_ctrl.vhdl:129:12  */
  always @*
    auto_data = n2892_q; // (isignal)
  initial
    auto_data = 32'b00000000000000000000000000000000;
  /* spi_flash_ctrl.vhdl:130:12  */
  always @*
    auto_cnt = n2893_q; // (isignal)
  initial
    auto_cnt = 6'b000000;
  /* spi_flash_ctrl.vhdl:131:12  */
  always @*
    auto_state = n2894_q; // (isignal)
  initial
    auto_state = 5'b00000;
  /* spi_flash_ctrl.vhdl:132:12  */
  assign auto_last_addr = n2895_q; // (signal)
  /* spi_flash_ctrl.vhdl:137:5  */
  spi_rxtx_4_1 spi_rxtx (
    .clk(clk),
    .rst(rst),
    .clk_div_i(cmd_clk_div),
    .cmd_valid_i(cmd_valid),
    .cmd_mode_i(cmd_mode),
    .cmd_clks_i(d_clks),
    .cmd_txd_i(d_tx),
    .sdat_i(sdat_i),
    .cmd_ready_o(spi_rxtx_cmd_ready_o),
    .d_rxd_o(spi_rxtx_d_rxd_o),
    .d_ack_o(spi_rxtx_d_ack_o),
    .bus_idle_o(spi_rxtx_bus_idle_o),
    .sck(spi_rxtx_sck),
    .sdat_o(spi_rxtx_sdat_o),
    .sdat_oe(spi_rxtx_sdat_oe));
  /* spi_flash_ctrl.vhdl:160:28  */
  assign n2044_o = wb_req[67];
  /* spi_flash_ctrl.vhdl:160:43  */
  assign n2045_o = wb_req[66];
  /* spi_flash_ctrl.vhdl:160:32  */
  assign n2046_o = n2044_o & n2045_o;
  /* spi_flash_ctrl.vhdl:161:30  */
  assign n2047_o = wb_valid & wb_sel_reg;
  /* spi_flash_ctrl.vhdl:162:30  */
  assign n2048_o = wb_valid & wb_sel_map;
  /* spi_flash_ctrl.vhdl:165:31  */
  assign n2049_o = wb_req[2:0];
  /* spi_flash_ctrl.vhdl:165:59  */
  assign n2050_o = wb_reg_valid ? n2049_o : 3'b111;
  /* spi_flash_ctrl.vhdl:168:37  */
  assign n2054_o = wb_reg == 3'b000;
  /* spi_flash_ctrl.vhdl:168:25  */
  assign n2055_o = n2054_o ? 1'b1 : 1'b0;
  /* spi_flash_ctrl.vhdl:181:32  */
  assign n2059_o = cmd_valid & cmd_ready;
  /* spi_flash_ctrl.vhdl:182:44  */
  assign n2060_o = wb_req[68];
  /* spi_flash_ctrl.vhdl:182:33  */
  assign n2061_o = ~n2060_o;
  /* spi_flash_ctrl.vhdl:183:13  */
  assign n2063_o = bus_idle ? 1'b0 : pending_read;
  /* spi_flash_ctrl.vhdl:181:13  */
  assign n2064_o = n2059_o ? n2061_o : n2063_o;
  assign n2068_o = ctrl_reg[1];
  /* spi_flash_ctrl.vhdl:193:73  */
  assign n2069_o = wb_req[68];
  /* spi_flash_ctrl.vhdl:193:62  */
  assign n2070_o = pending_read & n2069_o;
  /* spi_flash_ctrl.vhdl:193:44  */
  assign n2071_o = ~n2070_o;
  /* spi_flash_ctrl.vhdl:193:40  */
  assign n2072_o = wb_reg_dat_v & n2071_o;
  assign n2073_o = ctrl_reg[15:8];
  /* spi_flash_ctrl.vhdl:199:23  */
  assign n2075_o = wb_req[65:62];
  /* spi_flash_ctrl.vhdl:199:27  */
  assign n2077_o = n2075_o == 4'b0010;
  /* spi_flash_ctrl.vhdl:201:43  */
  assign n2078_o = wb_req[68];
  /* spi_flash_ctrl.vhdl:201:34  */
  assign n2080_o = {2'b10, n2078_o};
  /* spi_flash_ctrl.vhdl:203:26  */
  assign n2081_o = wb_req[65:62];
  /* spi_flash_ctrl.vhdl:203:30  */
  assign n2083_o = n2081_o == 4'b0100;
  /* spi_flash_ctrl.vhdl:205:43  */
  assign n2084_o = wb_req[68];
  /* spi_flash_ctrl.vhdl:205:34  */
  assign n2086_o = {2'b11, n2084_o};
  /* spi_flash_ctrl.vhdl:209:43  */
  assign n2087_o = wb_req[68];
  /* spi_flash_ctrl.vhdl:209:34  */
  assign n2089_o = {2'b01, n2087_o};
  /* spi_flash_ctrl.vhdl:203:13  */
  assign n2090_o = n2083_o ? n2086_o : n2089_o;
  /* spi_flash_ctrl.vhdl:203:13  */
  assign n2093_o = n2083_o ? 3'b001 : 3'b111;
  /* spi_flash_ctrl.vhdl:199:13  */
  assign n2094_o = n2077_o ? n2080_o : n2090_o;
  /* spi_flash_ctrl.vhdl:199:13  */
  assign n2096_o = n2077_o ? 3'b011 : n2093_o;
  /* spi_flash_ctrl.vhdl:212:37  */
  assign n2097_o = wb_req[37:30];
  assign n2098_o = ctrl_reg[1];
  /* spi_flash_ctrl.vhdl:213:27  */
  assign n2099_o = ~n2098_o;
  assign n2100_o = auto_cfg_reg[23:16];
  /* spi_flash_ctrl.vhdl:220:28  */
  assign n2102_o = ~auto_cs;
  /* spi_flash_ctrl.vhdl:191:9  */
  assign n2103_o = n2068_o ? n2099_o : n2102_o;
  /* spi_flash_ctrl.vhdl:191:9  */
  assign n2104_o = n2068_o ? n2072_o : auto_cmd_valid;
  /* spi_flash_ctrl.vhdl:191:9  */
  assign n2105_o = n2068_o ? n2073_o : n2100_o;
  /* spi_flash_ctrl.vhdl:191:9  */
  assign n2106_o = n2068_o ? n2094_o : auto_cmd_mode;
  /* spi_flash_ctrl.vhdl:191:9  */
  assign n2107_o = n2068_o ? n2096_o : auto_d_clks;
  /* spi_flash_ctrl.vhdl:191:9  */
  assign n2108_o = n2068_o ? n2097_o : auto_d_txd;
  /* spi_flash_ctrl.vhdl:247:27  */
  assign n2118_o = wb_rsp[33];
  /* spi_flash_ctrl.vhdl:247:50  */
  assign n2119_o = n2896_q[33];
  /* spi_flash_ctrl.vhdl:247:56  */
  assign n2120_o = ~n2119_o;
  /* spi_flash_ctrl.vhdl:247:39  */
  assign n2121_o = n2118_o & n2120_o;
  /* spi_flash_ctrl.vhdl:248:27  */
  assign n2122_o = n2023_o[66];
  /* spi_flash_ctrl.vhdl:247:62  */
  assign n2123_o = n2121_o & n2122_o;
  /* spi_flash_ctrl.vhdl:248:47  */
  assign n2124_o = n2023_o[67];
  /* spi_flash_ctrl.vhdl:248:37  */
  assign n2125_o = n2123_o & n2124_o;
  assign n2127_o = wb_rsp[33];
  /* spi_flash_ctrl.vhdl:247:17  */
  assign n2128_o = n2125_o ? 1'b1 : n2127_o;
  assign n2129_o = wb_rsp[32:0];
  /* spi_flash_ctrl.vhdl:247:17  */
  assign n2130_o = n2125_o ? n2023_o : wb_stash;
  /* spi_flash_ctrl.vhdl:254:27  */
  assign n2131_o = wb_rsp[33];
  /* spi_flash_ctrl.vhdl:254:33  */
  assign n2132_o = ~n2131_o;
  /* spi_flash_ctrl.vhdl:255:31  */
  assign n2133_o = n2896_q[33];
  /* spi_flash_ctrl.vhdl:261:34  */
  assign n2135_o = n2023_o[66];
  /* spi_flash_ctrl.vhdl:264:49  */
  assign n2136_o = n2023_o[66];
  /* spi_flash_ctrl.vhdl:265:49  */
  assign n2137_o = n2023_o[67];
  assign n2138_o = {n2137_o, n2136_o};
  assign n2139_o = n2023_o[65:0];
  assign n2140_o = wb_req[65:0];
  /* spi_flash_ctrl.vhdl:261:25  */
  assign n2141_o = n2135_o ? n2139_o : n2140_o;
  assign n2142_o = n2023_o[67:66];
  /* spi_flash_ctrl.vhdl:261:25  */
  assign n2143_o = n2135_o ? n2142_o : n2138_o;
  assign n2144_o = n2023_o[68];
  assign n2145_o = wb_req[68];
  /* spi_flash_ctrl.vhdl:261:25  */
  assign n2146_o = n2135_o ? n2144_o : n2145_o;
  /* spi_flash_ctrl.vhdl:254:17  */
  assign n2147_o = n2150_o ? 1'b0 : n2128_o;
  assign n2148_o = {n2146_o, n2143_o, n2141_o};
  /* spi_flash_ctrl.vhdl:255:21  */
  assign n2149_o = n2133_o ? wb_stash : n2148_o;
  /* spi_flash_ctrl.vhdl:254:17  */
  assign n2150_o = n2132_o & n2133_o;
  /* spi_flash_ctrl.vhdl:254:17  */
  assign n2151_o = n2132_o ? n2149_o : wb_req;
  assign n2152_o = {n2147_o, n2129_o};
  assign n2153_o = {1'b0, 1'b0};
  assign n2154_o = n2152_o[31:0];
  assign n2155_o = n2896_q[31:0];
  /* spi_flash_ctrl.vhdl:232:13  */
  assign n2156_o = rst ? n2155_o : n2154_o;
  assign n2157_o = n2152_o[33:32];
  /* spi_flash_ctrl.vhdl:232:13  */
  assign n2158_o = rst ? n2153_o : n2157_o;
  /* spi_flash_ctrl.vhdl:232:13  */
  assign n2159_o = rst ? wb_req : n2151_o;
  assign n2160_o = {1'b0, 1'b0, 1'b0, 4'b0000};
  assign n2161_o = n2130_o[61:0];
  assign n2162_o = wb_stash[61:0];
  /* spi_flash_ctrl.vhdl:232:13  */
  assign n2163_o = rst ? n2162_o : n2161_o;
  assign n2164_o = n2130_o[68:62];
  /* spi_flash_ctrl.vhdl:232:13  */
  assign n2165_o = rst ? n2160_o : n2164_o;
  assign n2166_o = {n2158_o, n2156_o};
  assign n2169_o = {n2165_o, n2163_o};
  /* spi_flash_ctrl.vhdl:277:29  */
  assign n2175_o = {8'b00000000, d_rx};
  /* spi_flash_ctrl.vhdl:277:36  */
  assign n2176_o = {n2175_o, d_rx};
  /* spi_flash_ctrl.vhdl:277:43  */
  assign n2177_o = {n2176_o, d_rx};
  /* spi_flash_ctrl.vhdl:284:29  */
  assign n2179_o = ~auto_ack;
  assign n2180_o = ctrl_reg[1];
  /* spi_flash_ctrl.vhdl:288:40  */
  assign n2182_o = wb_reg == 3'b000;
  /* spi_flash_ctrl.vhdl:288:29  */
  assign n2183_o = n2180_o & n2182_o;
  /* spi_flash_ctrl.vhdl:302:23  */
  assign n2184_o = wb_req[68];
  /* spi_flash_ctrl.vhdl:302:32  */
  assign n2185_o = n2184_o & pending_read;
  /* spi_flash_ctrl.vhdl:305:40  */
  assign n2187_o = wb_req[68];
  /* spi_flash_ctrl.vhdl:305:43  */
  assign n2188_o = n2187_o & cmd_ready;
  /* spi_flash_ctrl.vhdl:306:33  */
  assign n2189_o = ~cmd_ready;
  assign n2190_o = {n2189_o, n2188_o};
  assign n2191_o = n2190_o[0];
  /* spi_flash_ctrl.vhdl:302:13  */
  assign n2192_o = n2185_o ? 1'b0 : n2191_o;
  assign n2193_o = n2190_o[1];
  /* spi_flash_ctrl.vhdl:302:13  */
  assign n2194_o = n2185_o ? 1'b1 : n2193_o;
  /* spi_flash_ctrl.vhdl:317:27  */
  assign n2196_o = auto_state == 5'b00001;
  /* spi_flash_ctrl.vhdl:317:39  */
  assign n2197_o = n2196_o & bus_idle;
  assign n2216_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n2217_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n2218_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n2219_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n2220_o = {n2216_o, n2217_o, n2218_o, n2219_o};
  assign n2221_o = {n2220_o, ctrl_reg};
  /* spi_flash_ctrl.vhdl:322:17  */
  assign n2223_o = wb_reg == 3'b001;
  assign n2226_o = {1'b0, 1'b0, auto_cfg_reg};
  /* spi_flash_ctrl.vhdl:324:17  */
  assign n2228_o = wb_reg == 3'b010;
  assign n2229_o = {n2228_o, n2223_o};
  /* spi_flash_ctrl.vhdl:321:17  */
  always @*
    case (n2229_o)
      2'b10: n2230_o = n2226_o;
      2'b01: n2230_o = n2221_o;
      default: n2230_o = n2177_o;
    endcase
  assign n2232_o = {1'b0, 1'b1, n2230_o};
  assign n2233_o = n2232_o[32:0];
  assign n2234_o = {1'b0, n2177_o};
  /* spi_flash_ctrl.vhdl:317:13  */
  assign n2235_o = n2197_o ? n2233_o : n2234_o;
  assign n2236_o = n2232_o[33];
  /* spi_flash_ctrl.vhdl:317:13  */
  assign n2237_o = n2197_o ? n2236_o : 1'b1;
  assign n2238_o = {n2237_o, n2235_o};
  assign n2239_o = {1'b0, 1'b0, n2177_o};
  /* spi_flash_ctrl.vhdl:310:9  */
  assign n2240_o = wb_reg_valid ? n2238_o : n2239_o;
  assign n2241_o = {n2194_o, n2192_o};
  assign n2242_o = n2240_o[31:0];
  /* spi_flash_ctrl.vhdl:288:9  */
  assign n2243_o = n2183_o ? n2177_o : n2242_o;
  assign n2244_o = n2240_o[33:32];
  /* spi_flash_ctrl.vhdl:288:9  */
  assign n2245_o = n2183_o ? n2241_o : n2244_o;
  assign n2246_o = {n2245_o, n2243_o};
  assign n2247_o = {n2179_o, auto_ack, auto_data};
  assign n2249_o = ctrl_reg[1];
  /* spi_flash_ctrl.vhdl:341:26  */
  assign n2250_o = n2249_o & d_ack;
  assign n2252_o = n2247_o[32];
  assign n2253_o = n2246_o[32];
  /* spi_flash_ctrl.vhdl:281:9  */
  assign n2254_o = wb_map_valid ? n2252_o : n2253_o;
  /* spi_flash_ctrl.vhdl:341:9  */
  assign n2255_o = n2250_o ? 1'b1 : n2254_o;
  assign n2256_o = n2247_o[33];
  assign n2257_o = n2246_o[33];
  /* spi_flash_ctrl.vhdl:281:9  */
  assign n2258_o = wb_map_valid ? n2256_o : n2257_o;
  assign n2259_o = n2247_o[31:0];
  assign n2260_o = n2246_o[31:0];
  /* spi_flash_ctrl.vhdl:281:9  */
  assign n2261_o = wb_map_valid ? n2259_o : n2260_o;
  /* spi_flash_ctrl.vhdl:358:17  */
  assign n2265_o = auto_latch_adr ? auto_lad_next : auto_last_addr;
  /* spi_flash_ctrl.vhdl:351:13  */
  assign n2266_o = rst ? auto_data : auto_data_next;
  /* spi_flash_ctrl.vhdl:351:13  */
  assign n2267_o = rst ? auto_cnt : auto_cnt_next;
  /* spi_flash_ctrl.vhdl:351:13  */
  assign n2269_o = rst ? 5'b00000 : auto_next;
  /* spi_flash_ctrl.vhdl:351:13  */
  assign n2271_o = rst ? 32'b00000000000000000000000000000000 : n2265_o;
  /* spi_flash_ctrl.vhdl:396:34  */
  assign n2280_o = wb_req[27:0];
  /* spi_flash_ctrl.vhdl:396:22  */
  assign n2282_o = {2'b00, n2280_o};
  /* spi_flash_ctrl.vhdl:396:48  */
  assign n2284_o = {n2282_o, 2'b00};
  /* spi_flash_ctrl.vhdl:399:59  */
  assign n2286_o = n2284_o + 32'b00000000000000000000000000000100;
  /* spi_flash_ctrl.vhdl:402:29  */
  assign n2287_o = n2284_o == auto_last_addr;
  assign n2288_o = ctrl_reg[0];
  /* spi_flash_ctrl.vhdl:408:22  */
  assign n2289_o = rst | n2288_o;
  /* spi_flash_ctrl.vhdl:414:25  */
  assign n2290_o = {26'b0, auto_cnt};  //  uext
  /* spi_flash_ctrl.vhdl:414:25  */
  assign n2292_o = n2290_o != 32'b00000000000000000000000000000000;
  /* spi_flash_ctrl.vhdl:415:43  */
  assign n2293_o = {26'b0, auto_cnt};  //  uext
  /* spi_flash_ctrl.vhdl:415:43  */
  assign n2295_o = n2293_o - 32'b00000000000000000000000000000001;
  /* spi_flash_ctrl.vhdl:415:34  */
  assign n2296_o = n2295_o[5:0];  // trunc
  /* spi_flash_ctrl.vhdl:414:13  */
  assign n2297_o = n2292_o ? n2296_o : auto_cnt;
  /* spi_flash_ctrl.vhdl:419:28  */
  assign n2299_o = auto_state != 5'b00001;
  /* spi_flash_ctrl.vhdl:420:28  */
  assign n2301_o = auto_state != 5'b10011;
  /* spi_flash_ctrl.vhdl:419:41  */
  assign n2302_o = n2299_o & n2301_o;
  /* spi_flash_ctrl.vhdl:421:28  */
  assign n2304_o = auto_state != 5'b00000;
  /* spi_flash_ctrl.vhdl:420:45  */
  assign n2305_o = n2302_o & n2304_o;
  /* spi_flash_ctrl.vhdl:419:13  */
  assign n2308_o = n2305_o ? 1'b1 : 1'b0;
  /* spi_flash_ctrl.vhdl:427:13  */
  assign n2310_o = auto_state == 5'b00000;
  assign n2311_o = ctrl_reg[1];
  /* spi_flash_ctrl.vhdl:438:51  */
  assign n2312_o = ~n2311_o;
  /* spi_flash_ctrl.vhdl:438:39  */
  assign n2313_o = wb_map_valid & n2312_o;
  /* spi_flash_ctrl.vhdl:440:31  */
  assign n2314_o = wb_req[68];
  /* spi_flash_ctrl.vhdl:440:21  */
  assign n2316_o = n2314_o ? n2297_o : 6'b000001;
  /* spi_flash_ctrl.vhdl:440:21  */
  assign n2319_o = n2314_o ? 1'b1 : 1'b0;
  /* spi_flash_ctrl.vhdl:440:21  */
  assign n2321_o = n2314_o ? auto_state : 5'b00010;
  /* spi_flash_ctrl.vhdl:438:17  */
  assign n2322_o = n2313_o ? n2316_o : n2297_o;
  /* spi_flash_ctrl.vhdl:438:17  */
  assign n2324_o = n2313_o ? n2319_o : 1'b0;
  /* spi_flash_ctrl.vhdl:438:17  */
  assign n2325_o = n2313_o ? n2321_o : auto_state;
  /* spi_flash_ctrl.vhdl:436:13  */
  assign n2327_o = auto_state == 5'b00001;
  /* spi_flash_ctrl.vhdl:449:29  */
  assign n2328_o = {26'b0, auto_cnt};  //  uext
  /* spi_flash_ctrl.vhdl:449:29  */
  assign n2330_o = n2328_o == 32'b00000000000000000000000000000000;
  /* spi_flash_ctrl.vhdl:449:17  */
  assign n2332_o = n2330_o ? 5'b00011 : auto_state;
  /* spi_flash_ctrl.vhdl:448:13  */
  assign n2334_o = auto_state == 5'b00010;
  assign n2335_o = auto_cfg_reg[7:0];
  assign n2336_o = auto_cfg_reg[13];
  /* spi_flash_ctrl.vhdl:457:21  */
  assign n2339_o = n2336_o ? 5'b00111 : 5'b00110;
  /* spi_flash_ctrl.vhdl:456:17  */
  assign n2340_o = cmd_ready ? n2339_o : auto_state;
  /* spi_flash_ctrl.vhdl:453:13  */
  assign n2342_o = auto_state == 5'b00011;
  /* spi_flash_ctrl.vhdl:464:35  */
  assign n2343_o = n2284_o[31:24];
  /* spi_flash_ctrl.vhdl:466:17  */
  assign n2345_o = cmd_ready ? 5'b00110 : auto_state;
  /* spi_flash_ctrl.vhdl:463:13  */
  assign n2347_o = auto_state == 5'b00111;
  /* spi_flash_ctrl.vhdl:470:35  */
  assign n2348_o = n2284_o[23:16];
  /* spi_flash_ctrl.vhdl:472:17  */
  assign n2350_o = cmd_ready ? 5'b00101 : auto_state;
  /* spi_flash_ctrl.vhdl:469:13  */
  assign n2352_o = auto_state == 5'b00110;
  /* spi_flash_ctrl.vhdl:476:35  */
  assign n2353_o = n2284_o[15:8];
  /* spi_flash_ctrl.vhdl:478:17  */
  assign n2355_o = cmd_ready ? 5'b00100 : auto_state;
  /* spi_flash_ctrl.vhdl:475:13  */
  assign n2357_o = auto_state == 5'b00101;
  /* spi_flash_ctrl.vhdl:482:35  */
  assign n2358_o = n2284_o[7:0];
  assign n2360_o = auto_cfg_reg[10:8];
  /* spi_flash_ctrl.vhdl:485:41  */
  assign n2361_o = n2360_o == 3'b000;
  /* spi_flash_ctrl.vhdl:485:21  */
  assign n2364_o = n2361_o ? 5'b01001 : 5'b01000;
  /* spi_flash_ctrl.vhdl:484:17  */
  assign n2365_o = cmd_ready ? n2364_o : auto_state;
  /* spi_flash_ctrl.vhdl:481:13  */
  assign n2367_o = auto_state == 5'b00100;
  assign n2368_o = auto_cfg_reg[10:8];
  /* spi_flash_ctrl.vhdl:494:17  */
  assign n2370_o = cmd_ready ? 5'b01001 : auto_state;
  /* spi_flash_ctrl.vhdl:491:13  */
  assign n2372_o = auto_state == 5'b01000;
  assign n2373_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:499:48  */
  assign n2375_o = {n2373_o, 1'b0};
  assign n2382_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:371:21  */
  assign n2383_o = n2382_o == 2'b11;
  assign n2386_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:373:24  */
  assign n2387_o = n2386_o == 2'b10;
  /* spi_flash_ctrl.vhdl:373:13  */
  assign n2390_o = n2387_o ? 3'b011 : 3'b111;
  /* spi_flash_ctrl.vhdl:371:13  */
  assign n2391_o = n2383_o ? 3'b001 : n2390_o;
  /* spi_flash_ctrl.vhdl:501:17  */
  assign n2393_o = cmd_ready ? 5'b01101 : auto_state;
  /* spi_flash_ctrl.vhdl:497:13  */
  assign n2395_o = auto_state == 5'b01001;
  assign n2396_o = auto_data[7:0];
  /* spi_flash_ctrl.vhdl:505:17  */
  assign n2397_o = d_ack ? d_rx : n2396_o;
  /* spi_flash_ctrl.vhdl:505:17  */
  assign n2399_o = d_ack ? 5'b01010 : auto_state;
  /* spi_flash_ctrl.vhdl:504:13  */
  assign n2401_o = auto_state == 5'b01101;
  assign n2402_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:511:48  */
  assign n2404_o = {n2402_o, 1'b0};
  assign n2411_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:371:21  */
  assign n2412_o = n2411_o == 2'b11;
  assign n2415_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:373:24  */
  assign n2416_o = n2415_o == 2'b10;
  /* spi_flash_ctrl.vhdl:373:13  */
  assign n2419_o = n2416_o ? 3'b011 : 3'b111;
  /* spi_flash_ctrl.vhdl:371:13  */
  assign n2420_o = n2412_o ? 3'b001 : n2419_o;
  /* spi_flash_ctrl.vhdl:513:17  */
  assign n2422_o = cmd_ready ? 5'b01110 : auto_state;
  /* spi_flash_ctrl.vhdl:509:13  */
  assign n2424_o = auto_state == 5'b01010;
  assign n2425_o = auto_data[15:8];
  /* spi_flash_ctrl.vhdl:517:17  */
  assign n2426_o = d_ack ? d_rx : n2425_o;
  /* spi_flash_ctrl.vhdl:517:17  */
  assign n2428_o = d_ack ? 5'b01011 : auto_state;
  /* spi_flash_ctrl.vhdl:516:13  */
  assign n2430_o = auto_state == 5'b01110;
  assign n2431_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:523:48  */
  assign n2433_o = {n2431_o, 1'b0};
  assign n2440_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:371:21  */
  assign n2441_o = n2440_o == 2'b11;
  assign n2444_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:373:24  */
  assign n2445_o = n2444_o == 2'b10;
  /* spi_flash_ctrl.vhdl:373:13  */
  assign n2448_o = n2445_o ? 3'b011 : 3'b111;
  /* spi_flash_ctrl.vhdl:371:13  */
  assign n2449_o = n2441_o ? 3'b001 : n2448_o;
  /* spi_flash_ctrl.vhdl:525:17  */
  assign n2451_o = cmd_ready ? 5'b01111 : auto_state;
  /* spi_flash_ctrl.vhdl:521:13  */
  assign n2453_o = auto_state == 5'b01011;
  assign n2454_o = auto_data[23:16];
  /* spi_flash_ctrl.vhdl:529:17  */
  assign n2455_o = d_ack ? d_rx : n2454_o;
  /* spi_flash_ctrl.vhdl:529:17  */
  assign n2457_o = d_ack ? 5'b01100 : auto_state;
  /* spi_flash_ctrl.vhdl:528:13  */
  assign n2459_o = auto_state == 5'b01111;
  assign n2460_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:535:48  */
  assign n2462_o = {n2460_o, 1'b0};
  assign n2469_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:371:21  */
  assign n2470_o = n2469_o == 2'b11;
  assign n2473_o = auto_cfg_reg[12:11];
  /* spi_flash_ctrl.vhdl:373:24  */
  assign n2474_o = n2473_o == 2'b10;
  /* spi_flash_ctrl.vhdl:373:13  */
  assign n2477_o = n2474_o ? 3'b011 : 3'b111;
  /* spi_flash_ctrl.vhdl:371:13  */
  assign n2478_o = n2470_o ? 3'b001 : n2477_o;
  /* spi_flash_ctrl.vhdl:537:17  */
  assign n2480_o = cmd_ready ? 5'b10000 : auto_state;
  /* spi_flash_ctrl.vhdl:533:13  */
  assign n2482_o = auto_state == 5'b01100;
  assign n2483_o = auto_data[31:24];
  /* spi_flash_ctrl.vhdl:541:17  */
  assign n2484_o = d_ack ? d_rx : n2483_o;
  /* spi_flash_ctrl.vhdl:541:17  */
  assign n2486_o = d_ack ? 5'b10001 : auto_state;
  /* spi_flash_ctrl.vhdl:541:17  */
  assign n2489_o = d_ack ? 1'b1 : 1'b0;
  /* spi_flash_ctrl.vhdl:540:13  */
  assign n2491_o = auto_state == 5'b10000;
  assign n2492_o = auto_cfg_reg[29:24];
  /* spi_flash_ctrl.vhdl:546:13  */
  assign n2495_o = auto_state == 5'b10001;
  /* spi_flash_ctrl.vhdl:553:39  */
  assign n2496_o = wb_map_valid & n2287_o;
  /* spi_flash_ctrl.vhdl:553:66  */
  assign n2497_o = wb_req[68];
  /* spi_flash_ctrl.vhdl:553:69  */
  assign n2498_o = ~n2497_o;
  /* spi_flash_ctrl.vhdl:553:55  */
  assign n2499_o = n2496_o & n2498_o;
  /* spi_flash_ctrl.vhdl:555:42  */
  assign n2500_o = wb_map_valid | wb_reg_valid;
  /* spi_flash_ctrl.vhdl:555:76  */
  assign n2501_o = {26'b0, auto_cnt};  //  uext
  /* spi_flash_ctrl.vhdl:555:76  */
  assign n2503_o = n2501_o == 32'b00000000000000000000000000000000;
  /* spi_flash_ctrl.vhdl:555:64  */
  assign n2504_o = n2500_o | n2503_o;
  /* spi_flash_ctrl.vhdl:555:17  */
  assign n2506_o = n2504_o ? 6'b001010 : n2297_o;
  /* spi_flash_ctrl.vhdl:555:17  */
  assign n2508_o = n2504_o ? 5'b10011 : auto_state;
  /* spi_flash_ctrl.vhdl:553:17  */
  assign n2509_o = n2499_o ? n2297_o : n2506_o;
  /* spi_flash_ctrl.vhdl:553:17  */
  assign n2511_o = n2499_o ? 5'b01001 : n2508_o;
  /* spi_flash_ctrl.vhdl:550:13  */
  assign n2513_o = auto_state == 5'b10010;
  /* spi_flash_ctrl.vhdl:565:29  */
  assign n2514_o = {26'b0, auto_cnt};  //  uext
  /* spi_flash_ctrl.vhdl:565:29  */
  assign n2516_o = n2514_o == 32'b00000000000000000000000000000000;
  /* spi_flash_ctrl.vhdl:565:17  */
  assign n2518_o = n2516_o ? 5'b00001 : auto_state;
  /* spi_flash_ctrl.vhdl:564:13  */
  assign n2520_o = auto_state == 5'b10011;
  assign n2521_o = {n2520_o, n2513_o, n2495_o, n2491_o, n2482_o, n2459_o, n2453_o, n2430_o, n2424_o, n2401_o, n2395_o, n2372_o, n2367_o, n2357_o, n2352_o, n2347_o, n2342_o, n2334_o, n2327_o, n2310_o};
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2534_o = 1'b0;
      20'b01000000000000000000: n2534_o = 1'b0;
      20'b00100000000000000000: n2534_o = 1'b0;
      20'b00010000000000000000: n2534_o = 1'b0;
      20'b00001000000000000000: n2534_o = 1'b1;
      20'b00000100000000000000: n2534_o = 1'b0;
      20'b00000010000000000000: n2534_o = 1'b1;
      20'b00000001000000000000: n2534_o = 1'b0;
      20'b00000000100000000000: n2534_o = 1'b1;
      20'b00000000010000000000: n2534_o = 1'b0;
      20'b00000000001000000000: n2534_o = 1'b1;
      20'b00000000000100000000: n2534_o = 1'b1;
      20'b00000000000010000000: n2534_o = 1'b1;
      20'b00000000000001000000: n2534_o = 1'b1;
      20'b00000000000000100000: n2534_o = 1'b1;
      20'b00000000000000010000: n2534_o = 1'b1;
      20'b00000000000000001000: n2534_o = 1'b1;
      20'b00000000000000000100: n2534_o = 1'b0;
      20'b00000000000000000010: n2534_o = 1'b0;
      20'b00000000000000000001: n2534_o = 1'b0;
      default: n2534_o = 1'bX;
    endcase
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2537_o = 3'b001;
      20'b01000000000000000000: n2537_o = 3'b001;
      20'b00100000000000000000: n2537_o = 3'b001;
      20'b00010000000000000000: n2537_o = 3'b001;
      20'b00001000000000000000: n2537_o = n2462_o;
      20'b00000100000000000000: n2537_o = 3'b001;
      20'b00000010000000000000: n2537_o = n2433_o;
      20'b00000001000000000000: n2537_o = 3'b001;
      20'b00000000100000000000: n2537_o = n2404_o;
      20'b00000000010000000000: n2537_o = 3'b001;
      20'b00000000001000000000: n2537_o = n2375_o;
      20'b00000000000100000000: n2537_o = 3'b001;
      20'b00000000000010000000: n2537_o = 3'b001;
      20'b00000000000001000000: n2537_o = 3'b001;
      20'b00000000000000100000: n2537_o = 3'b001;
      20'b00000000000000010000: n2537_o = 3'b001;
      20'b00000000000000001000: n2537_o = 3'b001;
      20'b00000000000000000100: n2537_o = 3'b001;
      20'b00000000000000000010: n2537_o = 3'b001;
      20'b00000000000000000001: n2537_o = 3'b001;
      default: n2537_o = 3'bX;
    endcase
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2540_o = 8'b00000000;
      20'b01000000000000000000: n2540_o = 8'b00000000;
      20'b00100000000000000000: n2540_o = 8'b00000000;
      20'b00010000000000000000: n2540_o = 8'b00000000;
      20'b00001000000000000000: n2540_o = 8'b00000000;
      20'b00000100000000000000: n2540_o = 8'b00000000;
      20'b00000010000000000000: n2540_o = 8'b00000000;
      20'b00000001000000000000: n2540_o = 8'b00000000;
      20'b00000000100000000000: n2540_o = 8'b00000000;
      20'b00000000010000000000: n2540_o = 8'b00000000;
      20'b00000000001000000000: n2540_o = 8'b00000000;
      20'b00000000000100000000: n2540_o = 8'b00000000;
      20'b00000000000010000000: n2540_o = n2358_o;
      20'b00000000000001000000: n2540_o = n2353_o;
      20'b00000000000000100000: n2540_o = n2348_o;
      20'b00000000000000010000: n2540_o = n2343_o;
      20'b00000000000000001000: n2540_o = n2335_o;
      20'b00000000000000000100: n2540_o = 8'b00000000;
      20'b00000000000000000010: n2540_o = 8'b00000000;
      20'b00000000000000000001: n2540_o = 8'b00000000;
      default: n2540_o = 8'bX;
    endcase
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2543_o = 3'b111;
      20'b01000000000000000000: n2543_o = 3'b111;
      20'b00100000000000000000: n2543_o = 3'b111;
      20'b00010000000000000000: n2543_o = 3'b111;
      20'b00001000000000000000: n2543_o = n2478_o;
      20'b00000100000000000000: n2543_o = 3'b111;
      20'b00000010000000000000: n2543_o = n2449_o;
      20'b00000001000000000000: n2543_o = 3'b111;
      20'b00000000100000000000: n2543_o = n2420_o;
      20'b00000000010000000000: n2543_o = 3'b111;
      20'b00000000001000000000: n2543_o = n2391_o;
      20'b00000000000100000000: n2543_o = n2368_o;
      20'b00000000000010000000: n2543_o = 3'b111;
      20'b00000000000001000000: n2543_o = 3'b111;
      20'b00000000000000100000: n2543_o = 3'b111;
      20'b00000000000000010000: n2543_o = 3'b111;
      20'b00000000000000001000: n2543_o = 3'b111;
      20'b00000000000000000100: n2543_o = 3'b111;
      20'b00000000000000000010: n2543_o = 3'b111;
      20'b00000000000000000001: n2543_o = 3'b111;
      default: n2543_o = 3'bX;
    endcase
  assign n2544_o = auto_data[7:0];
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2546_o = n2544_o;
      20'b01000000000000000000: n2546_o = n2544_o;
      20'b00100000000000000000: n2546_o = n2544_o;
      20'b00010000000000000000: n2546_o = n2544_o;
      20'b00001000000000000000: n2546_o = n2544_o;
      20'b00000100000000000000: n2546_o = n2544_o;
      20'b00000010000000000000: n2546_o = n2544_o;
      20'b00000001000000000000: n2546_o = n2544_o;
      20'b00000000100000000000: n2546_o = n2544_o;
      20'b00000000010000000000: n2546_o = n2397_o;
      20'b00000000001000000000: n2546_o = n2544_o;
      20'b00000000000100000000: n2546_o = n2544_o;
      20'b00000000000010000000: n2546_o = n2544_o;
      20'b00000000000001000000: n2546_o = n2544_o;
      20'b00000000000000100000: n2546_o = n2544_o;
      20'b00000000000000010000: n2546_o = n2544_o;
      20'b00000000000000001000: n2546_o = n2544_o;
      20'b00000000000000000100: n2546_o = n2544_o;
      20'b00000000000000000010: n2546_o = n2544_o;
      20'b00000000000000000001: n2546_o = n2544_o;
      default: n2546_o = 8'bX;
    endcase
  assign n2547_o = auto_data[15:8];
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2549_o = n2547_o;
      20'b01000000000000000000: n2549_o = n2547_o;
      20'b00100000000000000000: n2549_o = n2547_o;
      20'b00010000000000000000: n2549_o = n2547_o;
      20'b00001000000000000000: n2549_o = n2547_o;
      20'b00000100000000000000: n2549_o = n2547_o;
      20'b00000010000000000000: n2549_o = n2547_o;
      20'b00000001000000000000: n2549_o = n2426_o;
      20'b00000000100000000000: n2549_o = n2547_o;
      20'b00000000010000000000: n2549_o = n2547_o;
      20'b00000000001000000000: n2549_o = n2547_o;
      20'b00000000000100000000: n2549_o = n2547_o;
      20'b00000000000010000000: n2549_o = n2547_o;
      20'b00000000000001000000: n2549_o = n2547_o;
      20'b00000000000000100000: n2549_o = n2547_o;
      20'b00000000000000010000: n2549_o = n2547_o;
      20'b00000000000000001000: n2549_o = n2547_o;
      20'b00000000000000000100: n2549_o = n2547_o;
      20'b00000000000000000010: n2549_o = n2547_o;
      20'b00000000000000000001: n2549_o = n2547_o;
      default: n2549_o = 8'bX;
    endcase
  assign n2550_o = auto_data[23:16];
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2552_o = n2550_o;
      20'b01000000000000000000: n2552_o = n2550_o;
      20'b00100000000000000000: n2552_o = n2550_o;
      20'b00010000000000000000: n2552_o = n2550_o;
      20'b00001000000000000000: n2552_o = n2550_o;
      20'b00000100000000000000: n2552_o = n2455_o;
      20'b00000010000000000000: n2552_o = n2550_o;
      20'b00000001000000000000: n2552_o = n2550_o;
      20'b00000000100000000000: n2552_o = n2550_o;
      20'b00000000010000000000: n2552_o = n2550_o;
      20'b00000000001000000000: n2552_o = n2550_o;
      20'b00000000000100000000: n2552_o = n2550_o;
      20'b00000000000010000000: n2552_o = n2550_o;
      20'b00000000000001000000: n2552_o = n2550_o;
      20'b00000000000000100000: n2552_o = n2550_o;
      20'b00000000000000010000: n2552_o = n2550_o;
      20'b00000000000000001000: n2552_o = n2550_o;
      20'b00000000000000000100: n2552_o = n2550_o;
      20'b00000000000000000010: n2552_o = n2550_o;
      20'b00000000000000000001: n2552_o = n2550_o;
      default: n2552_o = 8'bX;
    endcase
  assign n2553_o = auto_data[31:24];
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2555_o = n2553_o;
      20'b01000000000000000000: n2555_o = n2553_o;
      20'b00100000000000000000: n2555_o = n2553_o;
      20'b00010000000000000000: n2555_o = n2484_o;
      20'b00001000000000000000: n2555_o = n2553_o;
      20'b00000100000000000000: n2555_o = n2553_o;
      20'b00000010000000000000: n2555_o = n2553_o;
      20'b00000001000000000000: n2555_o = n2553_o;
      20'b00000000100000000000: n2555_o = n2553_o;
      20'b00000000010000000000: n2555_o = n2553_o;
      20'b00000000001000000000: n2555_o = n2553_o;
      20'b00000000000100000000: n2555_o = n2553_o;
      20'b00000000000010000000: n2555_o = n2553_o;
      20'b00000000000001000000: n2555_o = n2553_o;
      20'b00000000000000100000: n2555_o = n2553_o;
      20'b00000000000000010000: n2555_o = n2553_o;
      20'b00000000000000001000: n2555_o = n2553_o;
      20'b00000000000000000100: n2555_o = n2553_o;
      20'b00000000000000000010: n2555_o = n2553_o;
      20'b00000000000000000001: n2555_o = n2553_o;
      default: n2555_o = 8'bX;
    endcase
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2557_o = n2297_o;
      20'b01000000000000000000: n2557_o = n2509_o;
      20'b00100000000000000000: n2557_o = n2492_o;
      20'b00010000000000000000: n2557_o = n2297_o;
      20'b00001000000000000000: n2557_o = n2297_o;
      20'b00000100000000000000: n2557_o = n2297_o;
      20'b00000010000000000000: n2557_o = n2297_o;
      20'b00000001000000000000: n2557_o = n2297_o;
      20'b00000000100000000000: n2557_o = n2297_o;
      20'b00000000010000000000: n2557_o = n2297_o;
      20'b00000000001000000000: n2557_o = n2297_o;
      20'b00000000000100000000: n2557_o = n2297_o;
      20'b00000000000010000000: n2557_o = n2297_o;
      20'b00000000000001000000: n2557_o = n2297_o;
      20'b00000000000000100000: n2557_o = n2297_o;
      20'b00000000000000010000: n2557_o = n2297_o;
      20'b00000000000000001000: n2557_o = n2297_o;
      20'b00000000000000000100: n2557_o = n2297_o;
      20'b00000000000000000010: n2557_o = n2322_o;
      20'b00000000000000000001: n2557_o = n2297_o;
      default: n2557_o = 6'bX;
    endcase
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2561_o = 1'b0;
      20'b01000000000000000000: n2561_o = 1'b0;
      20'b00100000000000000000: n2561_o = 1'b1;
      20'b00010000000000000000: n2561_o = 1'b0;
      20'b00001000000000000000: n2561_o = 1'b0;
      20'b00000100000000000000: n2561_o = 1'b0;
      20'b00000010000000000000: n2561_o = 1'b0;
      20'b00000001000000000000: n2561_o = 1'b0;
      20'b00000000100000000000: n2561_o = 1'b0;
      20'b00000000010000000000: n2561_o = 1'b0;
      20'b00000000001000000000: n2561_o = 1'b0;
      20'b00000000000100000000: n2561_o = 1'b0;
      20'b00000000000010000000: n2561_o = 1'b0;
      20'b00000000000001000000: n2561_o = 1'b0;
      20'b00000000000000100000: n2561_o = 1'b0;
      20'b00000000000000010000: n2561_o = 1'b0;
      20'b00000000000000001000: n2561_o = 1'b0;
      20'b00000000000000000100: n2561_o = 1'b0;
      20'b00000000000000000010: n2561_o = n2324_o;
      20'b00000000000000000001: n2561_o = 1'b0;
      default: n2561_o = 1'bX;
    endcase
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2565_o = n2518_o;
      20'b01000000000000000000: n2565_o = n2511_o;
      20'b00100000000000000000: n2565_o = 5'b10010;
      20'b00010000000000000000: n2565_o = n2486_o;
      20'b00001000000000000000: n2565_o = n2480_o;
      20'b00000100000000000000: n2565_o = n2457_o;
      20'b00000010000000000000: n2565_o = n2451_o;
      20'b00000001000000000000: n2565_o = n2428_o;
      20'b00000000100000000000: n2565_o = n2422_o;
      20'b00000000010000000000: n2565_o = n2399_o;
      20'b00000000001000000000: n2565_o = n2393_o;
      20'b00000000000100000000: n2565_o = n2370_o;
      20'b00000000000010000000: n2565_o = n2365_o;
      20'b00000000000001000000: n2565_o = n2355_o;
      20'b00000000000000100000: n2565_o = n2350_o;
      20'b00000000000000010000: n2565_o = n2345_o;
      20'b00000000000000001000: n2565_o = n2340_o;
      20'b00000000000000000100: n2565_o = n2332_o;
      20'b00000000000000000010: n2565_o = n2325_o;
      20'b00000000000000000001: n2565_o = 5'b00001;
      default: n2565_o = 5'bX;
    endcase
  /* spi_flash_ctrl.vhdl:426:13  */
  always @*
    case (n2521_o)
      20'b10000000000000000000: n2568_o = 1'b0;
      20'b01000000000000000000: n2568_o = 1'b0;
      20'b00100000000000000000: n2568_o = 1'b0;
      20'b00010000000000000000: n2568_o = n2489_o;
      20'b00001000000000000000: n2568_o = 1'b0;
      20'b00000100000000000000: n2568_o = 1'b0;
      20'b00000010000000000000: n2568_o = 1'b0;
      20'b00000001000000000000: n2568_o = 1'b0;
      20'b00000000100000000000: n2568_o = 1'b0;
      20'b00000000010000000000: n2568_o = 1'b0;
      20'b00000000001000000000: n2568_o = 1'b0;
      20'b00000000000100000000: n2568_o = 1'b0;
      20'b00000000000010000000: n2568_o = 1'b0;
      20'b00000000000001000000: n2568_o = 1'b0;
      20'b00000000000000100000: n2568_o = 1'b0;
      20'b00000000000000010000: n2568_o = 1'b0;
      20'b00000000000000001000: n2568_o = 1'b0;
      20'b00000000000000000100: n2568_o = 1'b0;
      20'b00000000000000000010: n2568_o = 1'b0;
      20'b00000000000000000001: n2568_o = 1'b0;
      default: n2568_o = 1'bX;
    endcase
  /* spi_flash_ctrl.vhdl:408:9  */
  assign n2570_o = n2289_o ? 1'b0 : n2308_o;
  /* spi_flash_ctrl.vhdl:408:9  */
  assign n2573_o = n2289_o ? 1'b0 : n2534_o;
  /* spi_flash_ctrl.vhdl:408:9  */
  assign n2576_o = n2289_o ? 3'b001 : n2537_o;
  /* spi_flash_ctrl.vhdl:408:9  */
  assign n2579_o = n2289_o ? 8'b00000000 : n2540_o;
  /* spi_flash_ctrl.vhdl:408:9  */
  assign n2582_o = n2289_o ? 3'b111 : n2543_o;
  assign n2584_o = {n2555_o, n2552_o, n2549_o, n2546_o};
  /* spi_flash_ctrl.vhdl:408:9  */
  assign n2585_o = n2289_o ? auto_data : n2584_o;
  /* spi_flash_ctrl.vhdl:408:9  */
  assign n2587_o = n2289_o ? 6'b000000 : n2557_o;
  /* spi_flash_ctrl.vhdl:408:9  */
  assign n2589_o = n2289_o ? 1'b0 : n2561_o;
  /* spi_flash_ctrl.vhdl:408:9  */
  assign n2592_o = n2289_o ? 5'b00000 : n2565_o;
  /* spi_flash_ctrl.vhdl:408:9  */
  assign n2594_o = n2289_o ? 1'b0 : n2568_o;
  assign n2599_o = ctrl_reg[0];
  /* spi_flash_ctrl.vhdl:590:26  */
  assign n2600_o = rst | n2599_o;
  assign n2614_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n2615_o = ctrl_reg[3:0];
  /* spi_flash_ctrl.vhdl:590:13  */
  assign n2616_o = n2600_o ? n2614_o : n2615_o;
  assign n2617_o = ctrl_reg[15:8];
  /* spi_flash_ctrl.vhdl:590:13  */
  assign n2618_o = n2600_o ? 8'b00000100 : n2617_o;
  assign n2619_o = {6'b100000, 8'b00000100, 1'b0, 1'b0, 1'b0, 2'b00, 3'b000, 8'b00000011};
  /* spi_flash_ctrl.vhdl:590:13  */
  assign n2620_o = n2600_o ? n2619_o : auto_cfg_reg;
  /* spi_flash_ctrl.vhdl:612:46  */
  assign n2621_o = wb_req[68];
  /* spi_flash_ctrl.vhdl:612:35  */
  assign n2622_o = wb_reg_valid & n2621_o;
  /* spi_flash_ctrl.vhdl:612:70  */
  assign n2624_o = auto_state == 5'b00001;
  /* spi_flash_ctrl.vhdl:612:55  */
  assign n2625_o = n2622_o & n2624_o;
  /* spi_flash_ctrl.vhdl:612:82  */
  assign n2626_o = n2625_o & bus_idle;
  /* spi_flash_ctrl.vhdl:613:27  */
  assign n2628_o = wb_reg == 3'b001;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2637_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2638_o = wb_req[45];
  assign n2639_o = ctrl_reg[15];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2640_o = n2637_o ? n2638_o : n2639_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2642_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2643_o = wb_req[44];
  assign n2644_o = ctrl_reg[14];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2645_o = n2642_o ? n2643_o : n2644_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2647_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2648_o = wb_req[43];
  assign n2649_o = ctrl_reg[13];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2650_o = n2647_o ? n2648_o : n2649_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2652_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2653_o = wb_req[42];
  assign n2654_o = ctrl_reg[12];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2655_o = n2652_o ? n2653_o : n2654_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2657_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2658_o = wb_req[41];
  assign n2659_o = ctrl_reg[11];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2660_o = n2657_o ? n2658_o : n2659_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2662_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2663_o = wb_req[40];
  assign n2664_o = ctrl_reg[10];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2665_o = n2662_o ? n2663_o : n2664_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2667_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2668_o = wb_req[39];
  assign n2669_o = ctrl_reg[9];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2670_o = n2667_o ? n2668_o : n2669_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2672_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2673_o = wb_req[38];
  assign n2674_o = ctrl_reg[8];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2675_o = n2672_o ? n2673_o : n2674_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2677_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2678_o = wb_req[37];
  assign n2679_o = ctrl_reg[7];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2680_o = n2677_o ? n2678_o : n2679_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2682_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2683_o = wb_req[36];
  assign n2684_o = ctrl_reg[6];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2685_o = n2682_o ? n2683_o : n2684_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2687_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2688_o = wb_req[35];
  assign n2689_o = ctrl_reg[5];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2690_o = n2687_o ? n2688_o : n2689_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2692_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2693_o = wb_req[34];
  assign n2694_o = ctrl_reg[4];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2695_o = n2692_o ? n2693_o : n2694_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2697_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2698_o = wb_req[33];
  assign n2699_o = ctrl_reg[3];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2700_o = n2697_o ? n2698_o : n2699_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2702_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2703_o = wb_req[32];
  assign n2704_o = ctrl_reg[2];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2705_o = n2702_o ? n2703_o : n2704_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2707_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2708_o = wb_req[31];
  assign n2709_o = ctrl_reg[1];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2710_o = n2707_o ? n2708_o : n2709_o;
  assign n2711_o = ctrl_reg[0];
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2712_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2713_o = wb_req[30];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2714_o = n2712_o ? n2713_o : n2711_o;
  assign n2715_o = {n2640_o, n2645_o, n2650_o, n2655_o, n2660_o, n2665_o, n2670_o, n2675_o, n2680_o, n2685_o, n2690_o, n2695_o, n2700_o, n2705_o, n2710_o, n2714_o};
  assign n2716_o = ctrl_reg[7:4];
  assign n2717_o = {n2618_o, n2716_o, n2616_o};
  /* spi_flash_ctrl.vhdl:613:17  */
  assign n2718_o = n2628_o ? n2715_o : n2717_o;
  /* spi_flash_ctrl.vhdl:616:27  */
  assign n2720_o = wb_reg == 3'b010;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2729_o = wb_req[65];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2730_o = wb_req[59];
  assign n2731_o = auto_cfg_reg[29];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2732_o = n2729_o ? n2730_o : n2731_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2734_o = wb_req[65];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2735_o = wb_req[58];
  assign n2736_o = auto_cfg_reg[28];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2737_o = n2734_o ? n2735_o : n2736_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2739_o = wb_req[65];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2740_o = wb_req[57];
  assign n2741_o = auto_cfg_reg[27];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2742_o = n2739_o ? n2740_o : n2741_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2744_o = wb_req[65];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2745_o = wb_req[56];
  assign n2746_o = auto_cfg_reg[26];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2747_o = n2744_o ? n2745_o : n2746_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2749_o = wb_req[65];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2750_o = wb_req[55];
  assign n2751_o = auto_cfg_reg[25];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2752_o = n2749_o ? n2750_o : n2751_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2754_o = wb_req[65];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2755_o = wb_req[54];
  assign n2756_o = auto_cfg_reg[24];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2757_o = n2754_o ? n2755_o : n2756_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2759_o = wb_req[64];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2760_o = wb_req[53];
  assign n2761_o = auto_cfg_reg[23];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2762_o = n2759_o ? n2760_o : n2761_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2764_o = wb_req[64];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2765_o = wb_req[52];
  assign n2766_o = auto_cfg_reg[22];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2767_o = n2764_o ? n2765_o : n2766_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2769_o = wb_req[64];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2770_o = wb_req[51];
  assign n2771_o = auto_cfg_reg[21];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2772_o = n2769_o ? n2770_o : n2771_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2774_o = wb_req[64];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2775_o = wb_req[50];
  assign n2776_o = auto_cfg_reg[20];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2777_o = n2774_o ? n2775_o : n2776_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2779_o = wb_req[64];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2780_o = wb_req[49];
  assign n2781_o = auto_cfg_reg[19];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2782_o = n2779_o ? n2780_o : n2781_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2784_o = wb_req[64];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2785_o = wb_req[48];
  assign n2786_o = auto_cfg_reg[18];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2787_o = n2784_o ? n2785_o : n2786_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2789_o = wb_req[64];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2790_o = wb_req[47];
  assign n2791_o = auto_cfg_reg[17];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2792_o = n2789_o ? n2790_o : n2791_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2794_o = wb_req[64];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2795_o = wb_req[46];
  assign n2796_o = auto_cfg_reg[16];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2797_o = n2794_o ? n2795_o : n2796_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2799_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2800_o = wb_req[45];
  assign n2801_o = auto_cfg_reg[15];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2802_o = n2799_o ? n2800_o : n2801_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2804_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2805_o = wb_req[44];
  assign n2806_o = auto_cfg_reg[14];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2807_o = n2804_o ? n2805_o : n2806_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2809_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2810_o = wb_req[43];
  assign n2811_o = auto_cfg_reg[13];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2812_o = n2809_o ? n2810_o : n2811_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2814_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2815_o = wb_req[42];
  assign n2816_o = auto_cfg_reg[12];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2817_o = n2814_o ? n2815_o : n2816_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2819_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2820_o = wb_req[41];
  assign n2821_o = auto_cfg_reg[11];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2822_o = n2819_o ? n2820_o : n2821_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2824_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2825_o = wb_req[40];
  assign n2826_o = auto_cfg_reg[10];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2827_o = n2824_o ? n2825_o : n2826_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2829_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2830_o = wb_req[39];
  assign n2831_o = auto_cfg_reg[9];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2832_o = n2829_o ? n2830_o : n2831_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2834_o = wb_req[63];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2835_o = wb_req[38];
  assign n2836_o = auto_cfg_reg[8];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2837_o = n2834_o ? n2835_o : n2836_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2839_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2840_o = wb_req[37];
  assign n2841_o = auto_cfg_reg[7];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2842_o = n2839_o ? n2840_o : n2841_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2844_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2845_o = wb_req[36];
  assign n2846_o = auto_cfg_reg[6];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2847_o = n2844_o ? n2845_o : n2846_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2849_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2850_o = wb_req[35];
  assign n2851_o = auto_cfg_reg[5];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2852_o = n2849_o ? n2850_o : n2851_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2854_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2855_o = wb_req[34];
  assign n2856_o = auto_cfg_reg[4];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2857_o = n2854_o ? n2855_o : n2856_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2859_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2860_o = wb_req[33];
  assign n2861_o = auto_cfg_reg[3];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2862_o = n2859_o ? n2860_o : n2861_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2864_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2865_o = wb_req[32];
  assign n2866_o = auto_cfg_reg[2];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2867_o = n2864_o ? n2865_o : n2866_o;
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2869_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2870_o = wb_req[31];
  assign n2871_o = auto_cfg_reg[1];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2872_o = n2869_o ? n2870_o : n2871_o;
  assign n2873_o = auto_cfg_reg[0];
  /* spi_flash_ctrl.vhdl:581:25  */
  assign n2874_o = wb_req[62];
  /* spi_flash_ctrl.vhdl:582:34  */
  assign n2875_o = wb_req[30];
  /* spi_flash_ctrl.vhdl:581:17  */
  assign n2876_o = n2874_o ? n2875_o : n2873_o;
  assign n2877_o = {n2732_o, n2737_o, n2742_o, n2747_o, n2752_o, n2757_o, n2762_o, n2767_o, n2772_o, n2777_o, n2782_o, n2787_o, n2792_o, n2797_o, n2802_o, n2807_o, n2812_o, n2817_o, n2822_o, n2827_o, n2832_o, n2837_o, n2842_o, n2847_o, n2852_o, n2857_o, n2862_o, n2867_o, n2872_o, n2876_o};
  /* spi_flash_ctrl.vhdl:612:13  */
  assign n2878_o = n2882_o ? n2877_o : n2620_o;
  assign n2879_o = ctrl_reg[7:4];
  assign n2880_o = {n2618_o, n2879_o, n2616_o};
  /* spi_flash_ctrl.vhdl:612:13  */
  assign n2881_o = n2626_o ? n2718_o : n2880_o;
  /* spi_flash_ctrl.vhdl:612:13  */
  assign n2882_o = n2626_o & n2720_o;
  /* spi_flash_ctrl.vhdl:588:9  */
  always @(posedge clk)
    n2886_q <= n2881_o;
  initial
    n2886_q = 16'b0000000000000000;
  /* spi_flash_ctrl.vhdl:588:9  */
  always @(posedge clk)
    n2887_q <= n2878_o;
  initial
    n2887_q = 30'b000000000000000000000000000000;
  /* spi_flash_ctrl.vhdl:173:9  */
  always @(posedge clk)
    n2888_q <= n2064_o;
  /* spi_flash_ctrl.vhdl:231:9  */
  always @(posedge clk)
    n2889_q <= n2159_o;
  /* spi_flash_ctrl.vhdl:231:9  */
  always @(posedge clk)
    n2890_q <= n2169_o;
  /* spi_flash_ctrl.vhdl:231:9  */
  assign n2891_o = {n2258_o, n2255_o, n2261_o};
  /* spi_flash_ctrl.vhdl:350:9  */
  always @(posedge clk)
    n2892_q <= n2266_o;
  initial
    n2892_q = 32'b00000000000000000000000000000000;
  /* spi_flash_ctrl.vhdl:350:9  */
  always @(posedge clk)
    n2893_q <= n2267_o;
  initial
    n2893_q = 6'b000000;
  /* spi_flash_ctrl.vhdl:350:9  */
  always @(posedge clk)
    n2894_q <= n2269_o;
  initial
    n2894_q = 5'b00000;
  /* spi_flash_ctrl.vhdl:350:9  */
  always @(posedge clk)
    n2895_q <= n2271_o;
  /* spi_flash_ctrl.vhdl:231:9  */
  always @(posedge clk)
    n2896_q <= n2166_o;
endmodule

module syscon_100000000_4096_0_0_0_589433b711fb88bdee7cbb7d486960b51e4c8efd
  (input  clk,
   input  rst,
   input  [29:0] wishbone_in_adr,
   input  [31:0] wishbone_in_dat,
   input  [3:0] wishbone_in_sel,
   input  wishbone_in_cyc,
   input  wishbone_in_stb,
   input  wishbone_in_we,
   output [31:0] wishbone_out_dat,
   output wishbone_out_ack,
   output wishbone_out_stall,
   output dram_at_0,
   output core_reset,
   output soc_reset);
  wire [68:0] n1565_o;
  wire [31:0] n1567_o;
  wire n1568_o;
  wire n1569_o;
  wire [63:0] reg_out;
  wire [2:0] reg_ctrl;
  wire [63:0] reg_ctrl_out;
  wire [63:0] reg_info;
  wire [63:0] reg_braminfo;
  wire [63:0] reg_draminfo;
  wire [63:0] reg_dramiinfo;
  wire [63:0] reg_clkinfo;
  wire [63:0] reg_spiinfo;
  wire [63:0] reg_uart0info;
  wire [63:0] reg_uart1info;
  wire info_has_dram;
  wire info_has_bram;
  wire info_has_uart;
  wire info_has_spif;
  wire info_has_leth;
  wire info_has_lsdc;
  wire info_has_urt1;
  wire [39:0] info_clk;
  wire [31:0] info_fl_off;
  wire uinfo_16550;
  wire [31:0] uinfo_freq;
  wire [33:0] wb_rsp;
  wire n1575_o;
  wire n1576_o;
  wire n1577_o;
  wire n1578_o;
  wire n1581_o;
  wire n1585_o;
  wire n1589_o;
  wire n1593_o;
  wire n1597_o;
  wire n1601_o;
  wire n1605_o;
  wire [3:0] n1665_o;
  wire [3:0] n1666_o;
  wire [3:0] n1667_o;
  wire [3:0] n1668_o;
  wire [3:0] n1669_o;
  wire [3:0] n1670_o;
  wire [3:0] n1671_o;
  wire [3:0] n1672_o;
  wire [3:0] n1673_o;
  wire [3:0] n1674_o;
  wire [3:0] n1675_o;
  wire [3:0] n1676_o;
  wire [3:0] n1677_o;
  wire [3:0] n1678_o;
  wire [3:0] n1679_o;
  wire [3:0] n1680_o;
  wire [15:0] n1681_o;
  wire [15:0] n1682_o;
  wire [15:0] n1683_o;
  wire [15:0] n1684_o;
  wire [63:0] n1685_o;
  wire [63:0] n1689_o;
  wire [63:0] n1693_o;
  wire [3:0] n1719_o;
  wire [3:0] n1720_o;
  wire [3:0] n1721_o;
  wire [3:0] n1722_o;
  wire [3:0] n1723_o;
  wire [3:0] n1724_o;
  wire [15:0] n1725_o;
  wire [47:0] n1726_o;
  wire [63:0] n1727_o;
  wire [3:0] n1761_o;
  wire [3:0] n1762_o;
  wire [3:0] n1763_o;
  wire [3:0] n1764_o;
  wire [3:0] n1765_o;
  wire [3:0] n1766_o;
  wire [3:0] n1767_o;
  wire [3:0] n1768_o;
  wire [15:0] n1769_o;
  wire [15:0] n1770_o;
  wire [63:0] n1771_o;
  wire [3:0] n1833_o;
  wire [3:0] n1834_o;
  wire [3:0] n1835_o;
  wire [3:0] n1836_o;
  wire [3:0] n1837_o;
  wire [3:0] n1838_o;
  wire [3:0] n1839_o;
  wire [3:0] n1840_o;
  wire [3:0] n1841_o;
  wire [3:0] n1842_o;
  wire [3:0] n1843_o;
  wire [3:0] n1844_o;
  wire [3:0] n1845_o;
  wire [3:0] n1846_o;
  wire [3:0] n1847_o;
  wire [3:0] n1848_o;
  wire [15:0] n1849_o;
  wire [15:0] n1850_o;
  wire [15:0] n1851_o;
  wire [15:0] n1852_o;
  wire [63:0] n1853_o;
  wire n1856_o;
  wire [3:0] n1890_o;
  wire [3:0] n1891_o;
  wire [3:0] n1892_o;
  wire [3:0] n1893_o;
  wire [3:0] n1894_o;
  wire [3:0] n1895_o;
  wire [3:0] n1896_o;
  wire [3:0] n1897_o;
  wire [15:0] n1898_o;
  wire [15:0] n1899_o;
  wire [63:0] n1900_o;
  wire [3:0] n1933_o;
  wire [3:0] n1934_o;
  wire [3:0] n1935_o;
  wire [3:0] n1936_o;
  wire [3:0] n1937_o;
  wire [3:0] n1938_o;
  wire [3:0] n1939_o;
  wire [3:0] n1940_o;
  wire [15:0] n1941_o;
  wire [15:0] n1942_o;
  wire [63:0] n1943_o;
  wire n1944_o;
  wire n1945_o;
  wire n1946_o;
  wire [5:0] n1947_o;
  wire n1950_o;
  wire n1952_o;
  wire n1954_o;
  wire n1956_o;
  wire n1958_o;
  wire n1960_o;
  wire n1962_o;
  wire n1964_o;
  wire n1966_o;
  wire n1968_o;
  wire [9:0] n1970_o;
  reg [63:0] n1971_o;
  wire [31:0] n1972_o;
  wire n1973_o;
  wire [31:0] n1974_o;
  wire [31:0] n1975_o;
  wire n1983_o;
  wire n1984_o;
  wire n1985_o;
  wire n1986_o;
  wire n1987_o;
  wire [5:0] n1988_o;
  wire n1990_o;
  wire n1991_o;
  wire n1992_o;
  wire n1993_o;
  wire n1996_o;
  wire n1997_o;
  wire n1999_o;
  wire n2000_o;
  wire n2001_o;
  wire n2002_o;
  wire n2006_o;
  wire n2008_o;
  wire n2009_o;
  wire n2010_o;
  wire n2011_o;
  wire n2012_o;
  wire n2013_o;
  wire n2014_o;
  wire [2:0] n2015_o;
  wire [2:0] n2017_o;
  reg [2:0] n2020_q;
  wire [33:0] n2021_o;
  reg [33:0] n2022_q;
  assign wishbone_out_dat = n1567_o;
  assign wishbone_out_ack = n1568_o;
  assign wishbone_out_stall = n1569_o;
  assign dram_at_0 = n1575_o;
  assign core_reset = n1578_o;
  assign soc_reset = n1577_o;
  /* wishbone_arbiter.vhdl:38:39  */
  assign n1565_o = {wishbone_in_we, wishbone_in_stb, wishbone_in_cyc, wishbone_in_sel, wishbone_in_dat, wishbone_in_adr};
  assign n1567_o = n2022_q[31:0];
  assign n1568_o = n2022_q[32];
  assign n1569_o = n2022_q[33];
  /* syscon.vhdl:58:12  */
  assign reg_out = n1971_o; // (signal)
  /* syscon.vhdl:95:12  */
  assign reg_ctrl = n2020_q; // (signal)
  /* syscon.vhdl:96:12  */
  assign reg_ctrl_out = n1853_o; // (signal)
  /* syscon.vhdl:99:12  */
  assign reg_info = n1685_o; // (signal)
  /* syscon.vhdl:100:12  */
  assign reg_braminfo = 64'b0000000000000000000000000000000000000000000000000001000000000000; // (signal)
  /* syscon.vhdl:101:12  */
  assign reg_draminfo = n1689_o; // (signal)
  /* syscon.vhdl:102:12  */
  assign reg_dramiinfo = n1693_o; // (signal)
  /* syscon.vhdl:103:12  */
  assign reg_clkinfo = n1727_o; // (signal)
  /* syscon.vhdl:104:12  */
  assign reg_spiinfo = n1771_o; // (signal)
  /* syscon.vhdl:105:12  */
  assign reg_uart0info = n1900_o; // (signal)
  /* syscon.vhdl:106:12  */
  assign reg_uart1info = n1943_o; // (signal)
  /* syscon.vhdl:107:12  */
  assign info_has_dram = n1585_o; // (signal)
  /* syscon.vhdl:108:12  */
  assign info_has_bram = n1589_o; // (signal)
  /* syscon.vhdl:109:12  */
  assign info_has_uart = n1581_o; // (signal)
  /* syscon.vhdl:110:12  */
  assign info_has_spif = n1593_o; // (signal)
  /* syscon.vhdl:111:12  */
  assign info_has_leth = n1597_o; // (signal)
  /* syscon.vhdl:112:12  */
  assign info_has_lsdc = n1601_o; // (signal)
  /* syscon.vhdl:113:12  */
  assign info_has_urt1 = n1605_o; // (signal)
  /* syscon.vhdl:114:12  */
  assign info_clk = 40'b0000000000000101111101011110000100000000; // (signal)
  /* syscon.vhdl:115:12  */
  assign info_fl_off = 32'b00000000000000000000000000000000; // (signal)
  /* syscon.vhdl:116:12  */
  assign uinfo_16550 = n1856_o; // (signal)
  /* syscon.vhdl:117:12  */
  assign uinfo_freq = 32'b00000101111101011110000100000000; // (signal)
  /* syscon.vhdl:120:12  */
  assign wb_rsp = n2021_o; // (signal)
  /* syscon.vhdl:124:22  */
  assign n1575_o = 1'b0 ? 1'b1 : n1576_o;
  /* syscon.vhdl:124:54  */
  assign n1576_o = reg_ctrl[0];
  /* syscon.vhdl:125:26  */
  assign n1577_o = reg_ctrl[2];
  /* syscon.vhdl:126:27  */
  assign n1578_o = reg_ctrl[1];
  /* syscon.vhdl:129:26  */
  assign n1581_o = 1'b1 ? 1'b1 : 1'b0;
  /* syscon.vhdl:130:26  */
  assign n1585_o = 1'b1 ? 1'b1 : 1'b0;
  /* syscon.vhdl:131:26  */
  assign n1589_o = 1'b1 ? 1'b1 : 1'b0;
  /* syscon.vhdl:132:26  */
  assign n1593_o = 1'b1 ? 1'b1 : 1'b0;
  /* syscon.vhdl:133:26  */
  assign n1597_o = 1'b0 ? 1'b1 : 1'b0;
  /* syscon.vhdl:134:26  */
  assign n1601_o = 1'b0 ? 1'b1 : 1'b0;
  /* syscon.vhdl:135:26  */
  assign n1605_o = 1'b0 ? 1'b1 : 1'b0;
  assign n1665_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1666_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1667_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1668_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1669_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1670_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1671_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1672_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1673_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1674_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1675_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1676_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1677_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1678_o = {1'b0, 1'b0, 1'b0, info_has_lsdc};
  assign n1679_o = {1'b0, info_has_urt1, 1'b1, info_has_leth};
  assign n1680_o = {info_has_spif, info_has_bram, info_has_dram, info_has_uart};
  assign n1681_o = {n1665_o, n1666_o, n1667_o, n1668_o};
  assign n1682_o = {n1669_o, n1670_o, n1671_o, n1672_o};
  assign n1683_o = {n1673_o, n1674_o, n1675_o, n1676_o};
  assign n1684_o = {n1677_o, n1678_o, n1679_o, n1680_o};
  assign n1685_o = {n1681_o, n1682_o, n1683_o, n1684_o};
  /* syscon.vhdl:148:76  */
  assign n1689_o = 1'b1 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* syscon.vhdl:150:82  */
  assign n1693_o = 1'b1 ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  assign n1719_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1720_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1721_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1722_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1723_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1724_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1725_o = {n1719_o, n1720_o, n1721_o, n1722_o};
  assign n1726_o = {n1723_o, n1724_o, info_clk};
  assign n1727_o = {n1725_o, n1726_o};
  assign n1761_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1762_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1763_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1764_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1765_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1766_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1767_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1768_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1769_o = {n1761_o, n1762_o, n1763_o, n1764_o};
  assign n1770_o = {n1765_o, n1766_o, n1767_o, n1768_o};
  assign n1771_o = {n1769_o, n1770_o, info_fl_off};
  assign n1833_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1834_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1835_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1836_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1837_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1838_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1839_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1840_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1841_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1842_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1843_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1844_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1845_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1846_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1847_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1848_o = {1'b0, reg_ctrl};
  assign n1849_o = {n1833_o, n1834_o, n1835_o, n1836_o};
  assign n1850_o = {n1837_o, n1838_o, n1839_o, n1840_o};
  assign n1851_o = {n1841_o, n1842_o, n1843_o, n1844_o};
  assign n1852_o = {n1845_o, n1846_o, n1847_o, n1848_o};
  assign n1853_o = {n1849_o, n1850_o, n1851_o, n1852_o};
  /* syscon.vhdl:163:26  */
  assign n1856_o = 1'b1 ? 1'b1 : 1'b0;
  assign n1890_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1891_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1892_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1893_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1894_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1895_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1896_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1897_o = {1'b0, 1'b0, 1'b0, uinfo_16550};
  assign n1898_o = {n1890_o, n1891_o, n1892_o, n1893_o};
  assign n1899_o = {n1894_o, n1895_o, n1896_o, n1897_o};
  assign n1900_o = {n1898_o, n1899_o, uinfo_freq};
  assign n1933_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1934_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1935_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1936_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1937_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1938_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1939_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n1940_o = {1'b0, 1'b0, 1'b0, 1'b1};
  assign n1941_o = {n1933_o, n1934_o, n1935_o, n1936_o};
  assign n1942_o = {n1937_o, n1938_o, n1939_o, n1940_o};
  assign n1943_o = {n1941_o, n1942_o, uinfo_freq};
  /* syscon.vhdl:173:31  */
  assign n1944_o = n1565_o[66];
  /* syscon.vhdl:173:51  */
  assign n1945_o = n1565_o[67];
  /* syscon.vhdl:173:35  */
  assign n1946_o = n1944_o & n1945_o;
  /* syscon.vhdl:174:25  */
  assign n1947_o = n1565_o[6:1];
  /* syscon.vhdl:175:25  */
  assign n1950_o = n1947_o == 6'b000000;
  /* syscon.vhdl:176:25  */
  assign n1952_o = n1947_o == 6'b000001;
  /* syscon.vhdl:177:25  */
  assign n1954_o = n1947_o == 6'b000010;
  /* syscon.vhdl:178:25  */
  assign n1956_o = n1947_o == 6'b000011;
  /* syscon.vhdl:179:25  */
  assign n1958_o = n1947_o == 6'b000110;
  /* syscon.vhdl:180:25  */
  assign n1960_o = n1947_o == 6'b000100;
  /* syscon.vhdl:181:25  */
  assign n1962_o = n1947_o == 6'b000101;
  /* syscon.vhdl:182:25  */
  assign n1964_o = n1947_o == 6'b000111;
  /* syscon.vhdl:183:25  */
  assign n1966_o = n1947_o == 6'b001000;
  /* syscon.vhdl:184:25  */
  assign n1968_o = n1947_o == 6'b001001;
  assign n1970_o = {n1968_o, n1966_o, n1964_o, n1962_o, n1960_o, n1958_o, n1956_o, n1954_o, n1952_o, n1950_o};
  /* syscon.vhdl:174:5  */
  always @*
    case (n1970_o)
      10'b1000000000: n1971_o = reg_uart1info;
      10'b0100000000: n1971_o = reg_uart0info;
      10'b0010000000: n1971_o = reg_spiinfo;
      10'b0001000000: n1971_o = reg_ctrl_out;
      10'b0000100000: n1971_o = reg_clkinfo;
      10'b0000010000: n1971_o = reg_dramiinfo;
      10'b0000001000: n1971_o = reg_draminfo;
      10'b0000000100: n1971_o = reg_braminfo;
      10'b0000000010: n1971_o = reg_info;
      10'b0000000001: n1971_o = 64'b1111000000001101101010100101010100000000000000010000000000000001;
      default: n1971_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    endcase
  /* syscon.vhdl:186:28  */
  assign n1972_o = reg_out[63:32];
  /* syscon.vhdl:186:63  */
  assign n1973_o = n1565_o[0];
  /* syscon.vhdl:186:43  */
  assign n1974_o = n1973_o ? n1972_o : n1975_o;
  /* syscon.vhdl:187:26  */
  assign n1975_o = reg_out[31:0];
  /* syscon.vhdl:206:32  */
  assign n1983_o = n1565_o[66];
  /* syscon.vhdl:206:52  */
  assign n1984_o = n1565_o[67];
  /* syscon.vhdl:206:36  */
  assign n1985_o = n1983_o & n1984_o;
  /* syscon.vhdl:206:72  */
  assign n1986_o = n1565_o[68];
  /* syscon.vhdl:206:56  */
  assign n1987_o = n1985_o & n1986_o;
  /* syscon.vhdl:208:39  */
  assign n1988_o = n1565_o[6:1];
  /* syscon.vhdl:208:63  */
  assign n1990_o = n1988_o == 6'b000101;
  /* syscon.vhdl:209:40  */
  assign n1991_o = n1565_o[0];
  /* syscon.vhdl:209:44  */
  assign n1992_o = ~n1991_o;
  /* syscon.vhdl:208:78  */
  assign n1993_o = n1990_o & n1992_o;
  /* syscon.vhdl:206:17  */
  assign n1996_o = n1987_o & n1993_o;
  /* syscon.vhdl:216:28  */
  assign n1997_o = reg_ctrl[2];
  assign n1999_o = n1565_o[32];
  assign n2000_o = reg_ctrl[2];
  /* syscon.vhdl:206:17  */
  assign n2001_o = n1996_o ? n1999_o : n2000_o;
  /* syscon.vhdl:216:17  */
  assign n2002_o = n1997_o ? 1'b0 : n2001_o;
  /* syscon.vhdl:219:28  */
  assign n2006_o = reg_ctrl[1];
  assign n2008_o = n1565_o[31];
  assign n2009_o = reg_ctrl[1];
  /* syscon.vhdl:206:17  */
  assign n2010_o = n1996_o ? n2008_o : n2009_o;
  /* syscon.vhdl:219:17  */
  assign n2011_o = n2006_o ? 1'b0 : n2010_o;
  assign n2012_o = n1565_o[30];
  assign n2013_o = reg_ctrl[0];
  /* syscon.vhdl:206:17  */
  assign n2014_o = n1996_o ? n2012_o : n2013_o;
  assign n2015_o = {n2002_o, n2011_o, n2014_o};
  /* syscon.vhdl:203:13  */
  assign n2017_o = rst ? 3'b000 : n2015_o;
  /* syscon.vhdl:202:9  */
  always @(posedge clk)
    n2020_q <= n2017_o;
  /* syscon.vhdl:202:9  */
  assign n2021_o = {1'b0, n1946_o, n1974_o};
  /* syscon.vhdl:193:9  */
  always @(posedge clk)
    n2022_q <= wb_rsp;
endmodule

module wishbone_arbiter_4
  (input  clk,
   input  rst,
   input  [415:0] wb_masters_in,
   input  [63:0] wb_slave_in_dat,
   input  wb_slave_in_ack,
   input  wb_slave_in_stall,
   output [263:0] wb_masters_out,
   output [28:0] wb_slave_out_adr,
   output [63:0] wb_slave_out_dat,
   output [7:0] wb_slave_out_sel,
   output wb_slave_out_cyc,
   output wb_slave_out_stb,
   output wb_slave_out_we);
  wire [28:0] n1452_o;
  wire [63:0] n1453_o;
  wire [7:0] n1454_o;
  wire n1455_o;
  wire n1456_o;
  wire n1457_o;
  wire [65:0] n1458_o;
  wire [1:0] candidate;
  wire [1:0] selected;
  wire busy;
  wire [1:0] n1460_o;
  wire n1463_o;
  wire n1466_o;
  wire [1:0] n1467_o;
  wire [1:0] n1469_o;
  wire [63:0] n1472_o;
  wire n1473_o;
  wire [31:0] n1474_o;
  wire n1476_o;
  wire n1477_o;
  wire n1479_o;
  wire [31:0] n1480_o;
  wire n1482_o;
  wire n1483_o;
  wire [63:0] n1485_o;
  wire n1486_o;
  wire [31:0] n1487_o;
  wire n1489_o;
  wire n1490_o;
  wire n1492_o;
  wire [31:0] n1493_o;
  wire n1495_o;
  wire n1496_o;
  wire [63:0] n1498_o;
  wire n1499_o;
  wire [31:0] n1500_o;
  wire n1502_o;
  wire n1503_o;
  wire n1505_o;
  wire [31:0] n1506_o;
  wire n1508_o;
  wire n1509_o;
  wire [63:0] n1511_o;
  wire n1512_o;
  wire [31:0] n1513_o;
  wire n1515_o;
  wire n1516_o;
  wire n1518_o;
  wire [31:0] n1519_o;
  wire n1521_o;
  wire n1522_o;
  wire [103:0] n1526_o;
  wire n1527_o;
  wire [1:0] n1529_o;
  wire [103:0] n1530_o;
  wire n1531_o;
  wire [1:0] n1533_o;
  wire [103:0] n1534_o;
  wire n1535_o;
  wire [1:0] n1537_o;
  wire [103:0] n1538_o;
  wire n1539_o;
  wire [1:0] n1541_o;
  wire n1545_o;
  wire [1:0] n1546_o;
  wire [1:0] n1548_o;
  reg [1:0] n1551_q;
  wire [263:0] n1552_o;
  wire [103:0] n1553_o;
  wire [103:0] n1554_o;
  wire [103:0] n1555_o;
  wire [103:0] n1556_o;
  wire [1:0] n1557_o;
  reg [103:0] n1558_o;
  wire [103:0] n1559_o;
  wire [103:0] n1560_o;
  wire [103:0] n1561_o;
  wire [103:0] n1562_o;
  wire [1:0] n1563_o;
  reg [103:0] n1564_o;
  assign wb_masters_out = n1552_o;
  assign wb_slave_out_adr = n1452_o;
  assign wb_slave_out_dat = n1453_o;
  assign wb_slave_out_sel = n1454_o;
  assign wb_slave_out_cyc = n1455_o;
  assign wb_slave_out_stb = n1456_o;
  assign wb_slave_out_we = n1457_o;
  /* core.vhdl:489:29  */
  assign n1452_o = n1564_o[28:0];
  /* core.vhdl:487:28  */
  assign n1453_o = n1564_o[92:29];
  /* core.vhdl:482:27  */
  assign n1454_o = n1564_o[100:93];
  /* core.vhdl:481:25  */
  assign n1455_o = n1564_o[101];
  /* core.vhdl:480:26  */
  assign n1456_o = n1564_o[102];
  /* core.vhdl:479:24  */
  assign n1457_o = n1564_o[103];
  /* core.vhdl:476:25  */
  assign n1458_o = {wb_slave_in_stall, wb_slave_in_ack, wb_slave_in_dat};
  /* wishbone_arbiter.vhdl:25:12  */
  assign candidate = n1541_o; // (signal)
  /* wishbone_arbiter.vhdl:25:23  */
  assign selected = n1551_q; // (signal)
  /* wishbone_arbiter.vhdl:26:12  */
  assign busy = n1463_o; // (signal)
  /* wishbone_arbiter.vhdl:29:27  */
  assign n1460_o = 2'b11 - selected;
  /* wishbone_arbiter.vhdl:29:37  */
  assign n1463_o = n1558_o[101];
  /* wishbone_arbiter.vhdl:35:17  */
  assign n1466_o = ~busy;
  /* wishbone_arbiter.vhdl:35:9  */
  assign n1467_o = n1466_o ? candidate : selected;
  /* wishbone_arbiter.vhdl:38:39  */
  assign n1469_o = 2'b11 - n1467_o;
  /* wishbone_arbiter.vhdl:40:50  */
  assign n1472_o = n1458_o[63:0];
  /* wishbone_arbiter.vhdl:41:50  */
  assign n1473_o = n1458_o[64];
  /* wishbone_arbiter.vhdl:41:69  */
  assign n1474_o = {30'b0, n1467_o};  //  uext
  /* wishbone_arbiter.vhdl:41:69  */
  assign n1476_o = n1474_o == 32'b00000000000000000000000000000000;
  /* wishbone_arbiter.vhdl:41:54  */
  assign n1477_o = n1476_o ? n1473_o : 1'b0;
  /* wishbone_arbiter.vhdl:42:52  */
  assign n1479_o = n1458_o[65];
  /* wishbone_arbiter.vhdl:42:73  */
  assign n1480_o = {30'b0, n1467_o};  //  uext
  /* wishbone_arbiter.vhdl:42:73  */
  assign n1482_o = n1480_o == 32'b00000000000000000000000000000000;
  /* wishbone_arbiter.vhdl:42:58  */
  assign n1483_o = n1482_o ? n1479_o : 1'b1;
  /* wishbone_arbiter.vhdl:40:50  */
  assign n1485_o = n1458_o[63:0];
  /* wishbone_arbiter.vhdl:41:50  */
  assign n1486_o = n1458_o[64];
  /* wishbone_arbiter.vhdl:41:69  */
  assign n1487_o = {30'b0, n1467_o};  //  uext
  /* wishbone_arbiter.vhdl:41:69  */
  assign n1489_o = n1487_o == 32'b00000000000000000000000000000001;
  /* wishbone_arbiter.vhdl:41:54  */
  assign n1490_o = n1489_o ? n1486_o : 1'b0;
  /* wishbone_arbiter.vhdl:42:52  */
  assign n1492_o = n1458_o[65];
  /* wishbone_arbiter.vhdl:42:73  */
  assign n1493_o = {30'b0, n1467_o};  //  uext
  /* wishbone_arbiter.vhdl:42:73  */
  assign n1495_o = n1493_o == 32'b00000000000000000000000000000001;
  /* wishbone_arbiter.vhdl:42:58  */
  assign n1496_o = n1495_o ? n1492_o : 1'b1;
  /* wishbone_arbiter.vhdl:40:50  */
  assign n1498_o = n1458_o[63:0];
  /* wishbone_arbiter.vhdl:41:50  */
  assign n1499_o = n1458_o[64];
  /* wishbone_arbiter.vhdl:41:69  */
  assign n1500_o = {30'b0, n1467_o};  //  uext
  /* wishbone_arbiter.vhdl:41:69  */
  assign n1502_o = n1500_o == 32'b00000000000000000000000000000010;
  /* wishbone_arbiter.vhdl:41:54  */
  assign n1503_o = n1502_o ? n1499_o : 1'b0;
  /* wishbone_arbiter.vhdl:42:52  */
  assign n1505_o = n1458_o[65];
  /* wishbone_arbiter.vhdl:42:73  */
  assign n1506_o = {30'b0, n1467_o};  //  uext
  /* wishbone_arbiter.vhdl:42:73  */
  assign n1508_o = n1506_o == 32'b00000000000000000000000000000010;
  /* wishbone_arbiter.vhdl:42:58  */
  assign n1509_o = n1508_o ? n1505_o : 1'b1;
  /* wishbone_arbiter.vhdl:40:50  */
  assign n1511_o = n1458_o[63:0];
  /* wishbone_arbiter.vhdl:41:50  */
  assign n1512_o = n1458_o[64];
  /* wishbone_arbiter.vhdl:41:69  */
  assign n1513_o = {30'b0, n1467_o};  //  uext
  /* wishbone_arbiter.vhdl:41:69  */
  assign n1515_o = n1513_o == 32'b00000000000000000000000000000011;
  /* wishbone_arbiter.vhdl:41:54  */
  assign n1516_o = n1515_o ? n1512_o : 1'b0;
  /* wishbone_arbiter.vhdl:42:52  */
  assign n1518_o = n1458_o[65];
  /* wishbone_arbiter.vhdl:42:73  */
  assign n1519_o = {30'b0, n1467_o};  //  uext
  /* wishbone_arbiter.vhdl:42:73  */
  assign n1521_o = n1519_o == 32'b00000000000000000000000000000011;
  /* wishbone_arbiter.vhdl:42:58  */
  assign n1522_o = n1521_o ? n1518_o : 1'b1;
  /* wishbone_arbiter.vhdl:54:29  */
  assign n1526_o = wb_masters_in[103:0];
  /* wishbone_arbiter.vhdl:54:33  */
  assign n1527_o = n1526_o[101];
  /* wishbone_arbiter.vhdl:54:13  */
  assign n1529_o = n1527_o ? 2'b11 : selected;
  /* wishbone_arbiter.vhdl:54:29  */
  assign n1530_o = wb_masters_in[207:104];
  /* wishbone_arbiter.vhdl:54:33  */
  assign n1531_o = n1530_o[101];
  /* wishbone_arbiter.vhdl:54:13  */
  assign n1533_o = n1531_o ? 2'b10 : n1529_o;
  /* wishbone_arbiter.vhdl:54:29  */
  assign n1534_o = wb_masters_in[311:208];
  /* wishbone_arbiter.vhdl:54:33  */
  assign n1535_o = n1534_o[101];
  /* wishbone_arbiter.vhdl:54:13  */
  assign n1537_o = n1535_o ? 2'b01 : n1533_o;
  /* wishbone_arbiter.vhdl:54:29  */
  assign n1538_o = wb_masters_in[415:312];
  /* wishbone_arbiter.vhdl:54:33  */
  assign n1539_o = n1538_o[101];
  /* wishbone_arbiter.vhdl:54:13  */
  assign n1541_o = n1539_o ? 2'b00 : n1537_o;
  /* wishbone_arbiter.vhdl:65:24  */
  assign n1545_o = ~busy;
  /* wishbone_arbiter.vhdl:65:13  */
  assign n1546_o = n1545_o ? candidate : selected;
  /* wishbone_arbiter.vhdl:63:13  */
  assign n1548_o = rst ? 2'b00 : n1546_o;
  /* wishbone_arbiter.vhdl:62:9  */
  always @(posedge clk)
    n1551_q <= n1548_o;
  /* wishbone_arbiter.vhdl:62:9  */
  assign n1552_o = {n1483_o, n1477_o, n1472_o, n1496_o, n1490_o, n1485_o, n1509_o, n1503_o, n1498_o, n1522_o, n1516_o, n1511_o};
  /* wishbone_arbiter.vhdl:18:11  */
  assign n1553_o = wb_masters_in[103:0];
  /* wishbone_arbiter.vhdl:16:11  */
  assign n1554_o = wb_masters_in[207:104];
  assign n1555_o = wb_masters_in[311:208];
  /* wishbone_arbiter.vhdl:60:5  */
  assign n1556_o = wb_masters_in[415:312];
  /* wishbone_arbiter.vhdl:29:26  */
  assign n1557_o = n1460_o[1:0];
  /* wishbone_arbiter.vhdl:29:26  */
  always @*
    case (n1557_o)
      2'b00: n1558_o = n1553_o;
      2'b01: n1558_o = n1554_o;
      2'b10: n1558_o = n1555_o;
      2'b11: n1558_o = n1556_o;
    endcase
  /* wishbone_arbiter.vhdl:29:26  */
  assign n1559_o = wb_masters_in[103:0];
  /* wishbone_arbiter.vhdl:29:27  */
  assign n1560_o = wb_masters_in[207:104];
  /* core.vhdl:125:12  */
  assign n1561_o = wb_masters_in[311:208];
  /* wishbone_arbiter.vhdl:31:5  */
  assign n1562_o = wb_masters_in[415:312];
  /* wishbone_arbiter.vhdl:38:38  */
  assign n1563_o = n1469_o[1:0];
  /* wishbone_arbiter.vhdl:38:38  */
  always @*
    case (n1563_o)
      2'b00: n1564_o = n1559_o;
      2'b01: n1564_o = n1560_o;
      2'b10: n1564_o = n1561_o;
      2'b11: n1564_o = n1562_o;
    endcase
endmodule

module core_0_4_1_4_4_1_2_2_452bf2882a9b5f1c06340d5059c72dbd8af3bf8b
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  clk,
   input  rst,
   input  alt_reset,
   input  [63:0] wishbone_insn_in_dat,
   input  wishbone_insn_in_ack,
   input  wishbone_insn_in_stall,
   input  [63:0] wishbone_data_in_dat,
   input  wishbone_data_in_ack,
   input  wishbone_data_in_stall,
   input  [28:0] wb_snoop_in_adr,
   input  [63:0] wb_snoop_in_dat,
   input  [7:0] wb_snoop_in_sel,
   input  wb_snoop_in_cyc,
   input  wb_snoop_in_stb,
   input  wb_snoop_in_we,
   input  [3:0] dmi_addr,
   input  [63:0] dmi_din,
   input  dmi_req,
   input  dmi_wr,
   input  ext_irq,
   output [28:0] wishbone_insn_out_adr,
   output [63:0] wishbone_insn_out_dat,
   output [7:0] wishbone_insn_out_sel,
   output wishbone_insn_out_cyc,
   output wishbone_insn_out_stb,
   output wishbone_insn_out_we,
   output [28:0] wishbone_data_out_adr,
   output [63:0] wishbone_data_out_dat,
   output [7:0] wishbone_data_out_sel,
   output wishbone_data_out_cyc,
   output wishbone_data_out_stb,
   output wishbone_data_out_we,
   output [63:0] dmi_dout,
   output dmi_ack,
   output terminated_out);
  wire [65:0] n1004_o;
  wire [28:0] n1006_o;
  wire [63:0] n1007_o;
  wire [7:0] n1008_o;
  wire n1009_o;
  wire n1010_o;
  wire n1011_o;
  wire [65:0] n1012_o;
  wire [28:0] n1014_o;
  wire [63:0] n1015_o;
  wire [7:0] n1016_o;
  wire n1017_o;
  wire n1018_o;
  wire n1019_o;
  wire [103:0] n1020_o;
  wire [70:0] fetch1_to_icache;
  wire [134:0] writeback_to_fetch1;
  wire [101:0] icache_to_decode1;
  wire [130:0] mmu_to_icache;
  wire [164:0] decode1_to_decode2;
  wire [64:0] decode1_to_fetch1;
  wire [391:0] decode2_to_execute1;
  wire [191:0] register_file_to_decode2;
  wire [23:0] decode2_to_register_file;
  wire [71:0] writeback_to_register_file;
  wire decode2_to_cr_file;
  wire [36:0] cr_file_to_decode2;
  wire [46:0] writeback_to_cr_file;
  wire [353:0] execute1_to_writeback;
  wire [66:0] execute1_bypass;
  wire [34:0] execute1_cr_bypass;
  wire [389:0] execute1_to_loadstore1;
  wire [2:0] loadstore1_to_execute1;
  wire [175:0] loadstore1_to_writeback;
  wire [144:0] loadstore1_to_mmu;
  wire [70:0] mmu_to_loadstore1;
  wire [145:0] loadstore1_to_dcache;
  wire [67:0] dcache_to_loadstore1;
  wire [131:0] mmu_to_dcache;
  wire [66:0] dcache_to_mmu;
  wire [309:0] execute1_to_fpu;
  wire [1:0] fpu_to_execute1;
  wire [209:0] fpu_to_writeback;
  wire fetch1_stall_in;
  wire icache_stall_out;
  wire icache_stall_in;
  wire decode1_stall_in;
  wire decode1_busy;
  wire decode2_busy_in;
  wire decode2_stall_out;
  wire ex1_icache_inval;
  wire ex1_busy_out;
  wire dcache_stall_out;
  wire flush;
  wire decode1_flush;
  wire fetch1_flush;
  wire [2:0] complete;
  wire terminate;
  wire core_rst;
  wire do_interrupt;
  reg rst_fetch1;
  reg rst_icache;
  reg rst_dcache;
  reg rst_dec1;
  reg rst_dec2;
  reg rst_ex1;
  reg rst_fpu;
  reg rst_ls1;
  reg rst_wback;
  reg rst_dbg;
  wire alt_reset_d;
  wire sim_cr_dump;
  wire dbg_core_stop;
  wire dbg_core_rst;
  wire dbg_icache_rst;
  wire dbg_gpr_req;
  wire dbg_gpr_ack;
  wire [6:0] dbg_gpr_addr;
  wire [63:0] dbg_gpr_data;
  wire [63:0] msr;
  wire [1:0] icache_events;
  wire [2:0] loadstore_events;
  wire [4:0] dcache_events;
  wire [1:0] writeback_events;
  wire dbg_core_is_stopped;
  wire [255:0] log_data;
  wire [31:0] log_rd_addr;
  wire [31:0] log_wr_addr;
  wire [63:0] log_rd_data;
  wire n1035_o;
  wire fetch1_0_i_out_req;
  wire fetch1_0_i_out_virt_mode;
  wire fetch1_0_i_out_priv_mode;
  wire fetch1_0_i_out_big_endian;
  wire fetch1_0_i_out_stop_mark;
  wire fetch1_0_i_out_predicted;
  wire fetch1_0_i_out_pred_ntaken;
  wire [63:0] fetch1_0_i_out_nia;
  wire [42:0] fetch1_0_log_out;
  wire n1051_o;
  wire n1052_o;
  wire n1053_o;
  wire n1054_o;
  wire n1055_o;
  wire n1056_o;
  wire n1057_o;
  wire [63:0] n1058_o;
  wire [63:0] n1059_o;
  wire n1060_o;
  wire n1061_o;
  wire n1062_o;
  wire [63:0] n1063_o;
  wire [70:0] n1064_o;
  wire n1067_o;
  wire n1068_o;
  wire icache_0_i_out_valid;
  wire icache_0_i_out_stop_mark;
  wire icache_0_i_out_fetch_failed;
  wire [63:0] icache_0_i_out_nia;
  wire [31:0] icache_0_i_out_insn;
  wire icache_0_i_out_big_endian;
  wire icache_0_i_out_next_predicted;
  wire icache_0_i_out_next_pred_ntaken;
  wire icache_0_stall_out;
  wire [28:0] icache_0_wishbone_out_adr;
  wire [63:0] icache_0_wishbone_out_dat;
  wire [7:0] icache_0_wishbone_out_sel;
  wire icache_0_wishbone_out_cyc;
  wire icache_0_wishbone_out_stb;
  wire icache_0_wishbone_out_we;
  wire icache_0_events_icache_miss;
  wire icache_0_events_itlb_miss_resolved;
  wire [53:0] icache_0_log_out;
  wire n1069_o;
  wire n1070_o;
  wire n1071_o;
  wire n1072_o;
  wire n1073_o;
  wire n1074_o;
  wire n1075_o;
  wire [63:0] n1076_o;
  wire [101:0] n1077_o;
  wire n1079_o;
  wire n1080_o;
  wire n1081_o;
  wire [63:0] n1082_o;
  wire [63:0] n1083_o;
  wire n1085_o;
  wire [103:0] n1086_o;
  wire [63:0] n1088_o;
  wire n1089_o;
  wire n1090_o;
  wire [28:0] n1091_o;
  wire [63:0] n1092_o;
  wire [7:0] n1093_o;
  wire n1094_o;
  wire n1095_o;
  wire n1096_o;
  wire [1:0] n1097_o;
  wire decode1_0_busy_out;
  wire decode1_0_flush_out;
  wire decode1_0_f_out_redirect;
  wire [63:0] decode1_0_f_out_redirect_nia;
  wire decode1_0_d_out_valid;
  wire decode1_0_d_out_stop_mark;
  wire [63:0] decode1_0_d_out_nia;
  wire [31:0] decode1_0_d_out_insn;
  wire [6:0] decode1_0_d_out_ispr1;
  wire [6:0] decode1_0_d_out_ispr2;
  wire [6:0] decode1_0_d_out_ispro;
  wire [43:0] decode1_0_d_out_decode;
  wire decode1_0_d_out_br_pred;
  wire decode1_0_d_out_big_endian;
  wire [12:0] decode1_0_log_out;
  wire n1102_o;
  wire n1103_o;
  wire n1104_o;
  wire [63:0] n1105_o;
  wire [31:0] n1106_o;
  wire n1107_o;
  wire n1108_o;
  wire n1109_o;
  wire [64:0] n1110_o;
  wire [164:0] n1112_o;
  wire decode2_0_stall_out;
  wire decode2_0_stopped_out;
  wire decode2_0_e_out_valid;
  wire [1:0] decode2_0_e_out_unit;
  wire decode2_0_e_out_fac;
  wire [5:0] decode2_0_e_out_insn_type;
  wire [63:0] decode2_0_e_out_nia;
  wire [2:0] decode2_0_e_out_instr_tag;
  wire [6:0] decode2_0_e_out_write_reg;
  wire decode2_0_e_out_write_reg_enable;
  wire [6:0] decode2_0_e_out_read_reg1;
  wire [6:0] decode2_0_e_out_read_reg2;
  wire [63:0] decode2_0_e_out_read_data1;
  wire [63:0] decode2_0_e_out_read_data2;
  wire [63:0] decode2_0_e_out_read_data3;
  wire [31:0] decode2_0_e_out_cr;
  wire [4:0] decode2_0_e_out_xerc;
  wire decode2_0_e_out_lr;
  wire decode2_0_e_out_br_abs;
  wire decode2_0_e_out_rc;
  wire decode2_0_e_out_oe;
  wire decode2_0_e_out_invert_a;
  wire decode2_0_e_out_addm1;
  wire decode2_0_e_out_invert_out;
  wire [1:0] decode2_0_e_out_input_carry;
  wire decode2_0_e_out_output_carry;
  wire decode2_0_e_out_input_cr;
  wire decode2_0_e_out_output_cr;
  wire decode2_0_e_out_output_xer;
  wire decode2_0_e_out_is_32bit;
  wire decode2_0_e_out_is_signed;
  wire [31:0] decode2_0_e_out_insn;
  wire [3:0] decode2_0_e_out_data_len;
  wire decode2_0_e_out_byte_reverse;
  wire decode2_0_e_out_sign_extend;
  wire decode2_0_e_out_update;
  wire decode2_0_e_out_reserve;
  wire decode2_0_e_out_br_pred;
  wire [2:0] decode2_0_e_out_result_sel;
  wire [2:0] decode2_0_e_out_sub_select;
  wire decode2_0_e_out_repeat;
  wire decode2_0_e_out_second;
  wire decode2_0_r_out_read1_enable;
  wire [6:0] decode2_0_r_out_read1_reg;
  wire decode2_0_r_out_read2_enable;
  wire [6:0] decode2_0_r_out_read2_reg;
  wire decode2_0_r_out_read3_enable;
  wire [6:0] decode2_0_r_out_read3_reg;
  wire decode2_0_c_out_read;
  wire [9:0] decode2_0_log_out;
  wire [1:0] n1115_o;
  wire n1116_o;
  wire n1119_o;
  wire n1120_o;
  wire [63:0] n1121_o;
  wire [31:0] n1122_o;
  wire [6:0] n1123_o;
  wire [6:0] n1124_o;
  wire [6:0] n1125_o;
  wire [43:0] n1126_o;
  wire n1127_o;
  wire n1128_o;
  wire [391:0] n1129_o;
  wire [63:0] n1131_o;
  wire [63:0] n1132_o;
  wire [63:0] n1133_o;
  wire [23:0] n1134_o;
  wire [31:0] n1136_o;
  wire [4:0] n1137_o;
  wire [2:0] n1139_o;
  wire [63:0] n1140_o;
  wire [2:0] n1141_o;
  wire [31:0] n1142_o;
  wire [63:0] register_file_0_d_out_read1_data;
  wire [63:0] register_file_0_d_out_read2_data;
  wire [63:0] register_file_0_d_out_read3_data;
  wire register_file_0_dbg_gpr_ack;
  wire [63:0] register_file_0_dbg_gpr_data;
  wire register_file_0_sim_dump_done;
  wire [71:0] register_file_0_log_out;
  wire n1144_o;
  wire [6:0] n1145_o;
  wire n1146_o;
  wire [6:0] n1147_o;
  wire n1148_o;
  wire [6:0] n1149_o;
  wire [191:0] n1150_o;
  wire [6:0] n1152_o;
  wire [63:0] n1153_o;
  wire n1154_o;
  wire [31:0] cr_file_0_d_out_read_cr_data;
  wire [4:0] cr_file_0_d_out_read_xerc_data;
  wire [12:0] cr_file_0_log_out;
  wire n1159_o;
  wire [36:0] n1160_o;
  wire n1162_o;
  wire [7:0] n1163_o;
  wire [31:0] n1164_o;
  wire n1165_o;
  wire [4:0] n1166_o;
  wire execute1_0_busy_out;
  wire execute1_0_l_out_valid;
  wire [5:0] execute1_0_l_out_op;
  wire [63:0] execute1_0_l_out_nia;
  wire [31:0] execute1_0_l_out_insn;
  wire [2:0] execute1_0_l_out_instr_tag;
  wire [63:0] execute1_0_l_out_addr1;
  wire [63:0] execute1_0_l_out_addr2;
  wire [63:0] execute1_0_l_out_data;
  wire [6:0] execute1_0_l_out_write_reg;
  wire [3:0] execute1_0_l_out_length;
  wire execute1_0_l_out_ci;
  wire execute1_0_l_out_byte_reverse;
  wire execute1_0_l_out_sign_extend;
  wire execute1_0_l_out_update;
  wire [4:0] execute1_0_l_out_xerc;
  wire execute1_0_l_out_reserve;
  wire execute1_0_l_out_rc;
  wire execute1_0_l_out_virt_mode;
  wire execute1_0_l_out_priv_mode;
  wire execute1_0_l_out_mode_32bit;
  wire execute1_0_l_out_is_32bit;
  wire execute1_0_l_out_repeat;
  wire execute1_0_l_out_second;
  wire [63:0] execute1_0_l_out_msr;
  wire execute1_0_fp_out_valid;
  wire [5:0] execute1_0_fp_out_op;
  wire [63:0] execute1_0_fp_out_nia;
  wire [2:0] execute1_0_fp_out_itag;
  wire [31:0] execute1_0_fp_out_insn;
  wire execute1_0_fp_out_single;
  wire [1:0] execute1_0_fp_out_fe_mode;
  wire [63:0] execute1_0_fp_out_fra;
  wire [63:0] execute1_0_fp_out_frb;
  wire [63:0] execute1_0_fp_out_frc;
  wire [6:0] execute1_0_fp_out_frt;
  wire execute1_0_fp_out_rc;
  wire execute1_0_fp_out_out_cr;
  wire execute1_0_e_out_valid;
  wire [2:0] execute1_0_e_out_instr_tag;
  wire execute1_0_e_out_rc;
  wire execute1_0_e_out_mode_32bit;
  wire execute1_0_e_out_write_enable;
  wire [6:0] execute1_0_e_out_write_reg;
  wire [63:0] execute1_0_e_out_write_data;
  wire execute1_0_e_out_write_cr_enable;
  wire [7:0] execute1_0_e_out_write_cr_mask;
  wire [31:0] execute1_0_e_out_write_cr_data;
  wire execute1_0_e_out_write_xerc_enable;
  wire [4:0] execute1_0_e_out_xerc;
  wire execute1_0_e_out_interrupt;
  wire [11:0] execute1_0_e_out_intr_vec;
  wire execute1_0_e_out_redirect;
  wire [3:0] execute1_0_e_out_redir_mode;
  wire [63:0] execute1_0_e_out_last_nia;
  wire [63:0] execute1_0_e_out_br_offset;
  wire execute1_0_e_out_br_last;
  wire execute1_0_e_out_br_taken;
  wire execute1_0_e_out_abs_br;
  wire [15:0] execute1_0_e_out_srr1;
  wire [63:0] execute1_0_e_out_msr;
  wire [2:0] execute1_0_bypass_data_tag;
  wire [63:0] execute1_0_bypass_data_data;
  wire [2:0] execute1_0_bypass_cr_data_tag;
  wire [31:0] execute1_0_bypass_cr_data_data;
  wire [63:0] execute1_0_dbg_msr_out;
  wire execute1_0_icache_inval;
  wire execute1_0_terminate_out;
  wire [14:0] execute1_0_log_out;
  wire [31:0] execute1_0_log_rd_addr;
  wire n1169_o;
  wire [1:0] n1170_o;
  wire n1171_o;
  wire [5:0] n1172_o;
  wire [63:0] n1173_o;
  wire [2:0] n1174_o;
  wire [6:0] n1175_o;
  wire n1176_o;
  wire [6:0] n1177_o;
  wire [6:0] n1178_o;
  wire [63:0] n1179_o;
  wire [63:0] n1180_o;
  wire [63:0] n1181_o;
  wire [31:0] n1182_o;
  wire [4:0] n1183_o;
  wire n1184_o;
  wire n1185_o;
  wire n1186_o;
  wire n1187_o;
  wire n1188_o;
  wire n1189_o;
  wire n1190_o;
  wire [1:0] n1191_o;
  wire n1192_o;
  wire n1193_o;
  wire n1194_o;
  wire n1195_o;
  wire n1196_o;
  wire n1197_o;
  wire [31:0] n1198_o;
  wire [3:0] n1199_o;
  wire n1200_o;
  wire n1201_o;
  wire n1202_o;
  wire n1203_o;
  wire n1204_o;
  wire [2:0] n1205_o;
  wire [2:0] n1206_o;
  wire n1207_o;
  wire n1208_o;
  wire n1209_o;
  wire n1210_o;
  wire n1211_o;
  wire n1212_o;
  wire n1213_o;
  wire [389:0] n1214_o;
  wire [309:0] n1216_o;
  wire [353:0] n1218_o;
  wire [66:0] n1220_o;
  wire [34:0] n1222_o;
  wire n1227_o;
  wire n1228_o;
  wire n1229_o;
  wire n1230_o;
  wire n1231_o;
  wire n1232_o;
  wire n1233_o;
  wire n1234_o;
  wire n1235_o;
  wire n1236_o;
  wire n1237_o;
  wire n1238_o;
  wire with_fpu_fpu_0_e_out_busy;
  wire with_fpu_fpu_0_e_out_exception;
  wire with_fpu_fpu_0_w_out_valid;
  wire with_fpu_fpu_0_w_out_interrupt;
  wire [2:0] with_fpu_fpu_0_w_out_instr_tag;
  wire with_fpu_fpu_0_w_out_write_enable;
  wire [6:0] with_fpu_fpu_0_w_out_write_reg;
  wire [63:0] with_fpu_fpu_0_w_out_write_data;
  wire with_fpu_fpu_0_w_out_write_cr_enable;
  wire [7:0] with_fpu_fpu_0_w_out_write_cr_mask;
  wire [31:0] with_fpu_fpu_0_w_out_write_cr_data;
  wire [11:0] with_fpu_fpu_0_w_out_intr_vec;
  wire [63:0] with_fpu_fpu_0_w_out_srr0;
  wire [15:0] with_fpu_fpu_0_w_out_srr1;
  wire n1241_o;
  wire [5:0] n1242_o;
  wire [63:0] n1243_o;
  wire [2:0] n1244_o;
  wire [31:0] n1245_o;
  wire n1246_o;
  wire [1:0] n1247_o;
  wire [63:0] n1248_o;
  wire [63:0] n1249_o;
  wire [63:0] n1250_o;
  wire [6:0] n1251_o;
  wire n1252_o;
  wire n1253_o;
  wire [1:0] n1254_o;
  wire [209:0] n1256_o;
  wire loadstore1_0_e_out_busy;
  wire loadstore1_0_e_out_in_progress;
  wire loadstore1_0_e_out_interrupt;
  wire loadstore1_0_l_out_valid;
  wire [2:0] loadstore1_0_l_out_instr_tag;
  wire loadstore1_0_l_out_write_enable;
  wire [6:0] loadstore1_0_l_out_write_reg;
  wire [63:0] loadstore1_0_l_out_write_data;
  wire [4:0] loadstore1_0_l_out_xerc;
  wire loadstore1_0_l_out_rc;
  wire loadstore1_0_l_out_store_done;
  wire loadstore1_0_l_out_interrupt;
  wire [11:0] loadstore1_0_l_out_intr_vec;
  wire [63:0] loadstore1_0_l_out_srr0;
  wire [15:0] loadstore1_0_l_out_srr1;
  wire loadstore1_0_d_out_valid;
  wire loadstore1_0_d_out_hold;
  wire loadstore1_0_d_out_load;
  wire loadstore1_0_d_out_dcbz;
  wire loadstore1_0_d_out_nc;
  wire loadstore1_0_d_out_reserve;
  wire loadstore1_0_d_out_atomic;
  wire loadstore1_0_d_out_atomic_last;
  wire loadstore1_0_d_out_virt_mode;
  wire loadstore1_0_d_out_priv_mode;
  wire [63:0] loadstore1_0_d_out_addr;
  wire [63:0] loadstore1_0_d_out_data;
  wire [7:0] loadstore1_0_d_out_byte_sel;
  wire loadstore1_0_m_out_valid;
  wire loadstore1_0_m_out_tlbie;
  wire loadstore1_0_m_out_slbia;
  wire loadstore1_0_m_out_mtspr;
  wire loadstore1_0_m_out_iside;
  wire loadstore1_0_m_out_load;
  wire loadstore1_0_m_out_priv;
  wire [9:0] loadstore1_0_m_out_sprn;
  wire [63:0] loadstore1_0_m_out_addr;
  wire [63:0] loadstore1_0_m_out_rs;
  wire loadstore1_0_events_load_complete;
  wire loadstore1_0_events_store_complete;
  wire loadstore1_0_events_itlb_miss;
  wire [9:0] loadstore1_0_log_out;
  wire n1258_o;
  wire [5:0] n1259_o;
  wire [63:0] n1260_o;
  wire [31:0] n1261_o;
  wire [2:0] n1262_o;
  wire [63:0] n1263_o;
  wire [63:0] n1264_o;
  wire [63:0] n1265_o;
  wire [6:0] n1266_o;
  wire [3:0] n1267_o;
  wire n1268_o;
  wire n1269_o;
  wire n1270_o;
  wire n1271_o;
  wire [4:0] n1272_o;
  wire n1273_o;
  wire n1274_o;
  wire n1275_o;
  wire n1276_o;
  wire n1277_o;
  wire n1278_o;
  wire n1279_o;
  wire n1280_o;
  wire [63:0] n1281_o;
  wire [2:0] n1282_o;
  wire [175:0] n1284_o;
  wire [145:0] n1286_o;
  wire n1288_o;
  wire [63:0] n1289_o;
  wire n1290_o;
  wire n1291_o;
  wire n1292_o;
  wire [144:0] n1293_o;
  wire n1295_o;
  wire n1296_o;
  wire n1297_o;
  wire n1298_o;
  wire n1299_o;
  wire n1300_o;
  wire n1301_o;
  wire [63:0] n1302_o;
  wire [2:0] n1303_o;
  wire mmu_0_l_out_done;
  wire mmu_0_l_out_err;
  wire mmu_0_l_out_invalid;
  wire mmu_0_l_out_badtree;
  wire mmu_0_l_out_segerr;
  wire mmu_0_l_out_perm_error;
  wire mmu_0_l_out_rc_error;
  wire [63:0] mmu_0_l_out_sprval;
  wire mmu_0_d_out_valid;
  wire mmu_0_d_out_tlbie;
  wire mmu_0_d_out_doall;
  wire mmu_0_d_out_tlbld;
  wire [63:0] mmu_0_d_out_addr;
  wire [63:0] mmu_0_d_out_pte;
  wire mmu_0_i_out_tlbld;
  wire mmu_0_i_out_tlbie;
  wire mmu_0_i_out_doall;
  wire [63:0] mmu_0_i_out_addr;
  wire [63:0] mmu_0_i_out_pte;
  wire n1306_o;
  wire n1307_o;
  wire n1308_o;
  wire n1309_o;
  wire n1310_o;
  wire n1311_o;
  wire n1312_o;
  wire [9:0] n1313_o;
  wire [63:0] n1314_o;
  wire [63:0] n1315_o;
  wire [70:0] n1316_o;
  wire [131:0] n1318_o;
  wire n1320_o;
  wire n1321_o;
  wire n1322_o;
  wire [63:0] n1323_o;
  wire [130:0] n1324_o;
  wire dcache_0_d_out_valid;
  wire [63:0] dcache_0_d_out_data;
  wire dcache_0_d_out_store_done;
  wire dcache_0_d_out_error;
  wire dcache_0_d_out_cache_paradox;
  wire dcache_0_m_out_stall;
  wire dcache_0_m_out_done;
  wire dcache_0_m_out_err;
  wire [63:0] dcache_0_m_out_data;
  wire dcache_0_stall_out;
  wire [28:0] dcache_0_wishbone_out_adr;
  wire [63:0] dcache_0_wishbone_out_dat;
  wire [7:0] dcache_0_wishbone_out_sel;
  wire dcache_0_wishbone_out_cyc;
  wire dcache_0_wishbone_out_stb;
  wire dcache_0_wishbone_out_we;
  wire dcache_0_events_load_miss;
  wire dcache_0_events_store_miss;
  wire dcache_0_events_dcache_refill;
  wire dcache_0_events_dtlb_miss;
  wire dcache_0_events_dtlb_miss_resolved;
  wire [19:0] dcache_0_log_out;
  wire n1326_o;
  wire n1327_o;
  wire n1328_o;
  wire n1329_o;
  wire n1330_o;
  wire n1331_o;
  wire n1332_o;
  wire n1333_o;
  wire n1334_o;
  wire n1335_o;
  wire [63:0] n1336_o;
  wire [63:0] n1337_o;
  wire [7:0] n1338_o;
  wire [67:0] n1339_o;
  wire n1341_o;
  wire n1342_o;
  wire n1343_o;
  wire n1344_o;
  wire [63:0] n1345_o;
  wire [63:0] n1346_o;
  wire [66:0] n1347_o;
  wire [28:0] n1349_o;
  wire [63:0] n1350_o;
  wire [7:0] n1351_o;
  wire n1352_o;
  wire n1353_o;
  wire n1354_o;
  wire [103:0] n1356_o;
  wire [63:0] n1358_o;
  wire n1359_o;
  wire n1360_o;
  wire [4:0] n1361_o;
  wire [6:0] writeback_0_w_out_write_reg;
  wire [63:0] writeback_0_w_out_write_data;
  wire writeback_0_w_out_write_enable;
  wire writeback_0_c_out_write_cr_enable;
  wire [7:0] writeback_0_c_out_write_cr_mask;
  wire [31:0] writeback_0_c_out_write_cr_data;
  wire writeback_0_c_out_write_xerc_enable;
  wire [4:0] writeback_0_c_out_write_xerc_data;
  wire writeback_0_f_out_redirect;
  wire writeback_0_f_out_virt_mode;
  wire writeback_0_f_out_priv_mode;
  wire writeback_0_f_out_big_endian;
  wire writeback_0_f_out_mode_32bit;
  wire [63:0] writeback_0_f_out_redirect_nia;
  wire [63:0] writeback_0_f_out_br_nia;
  wire writeback_0_f_out_br_last;
  wire writeback_0_f_out_br_taken;
  wire writeback_0_events_instr_complete;
  wire writeback_0_events_fp_complete;
  wire writeback_0_flush_out;
  wire writeback_0_interrupt_out;
  wire [1:0] writeback_0_complete_out_tag;
  wire writeback_0_complete_out_valid;
  wire n1364_o;
  wire [2:0] n1365_o;
  wire n1366_o;
  wire n1367_o;
  wire n1368_o;
  wire [6:0] n1369_o;
  wire [63:0] n1370_o;
  wire n1371_o;
  wire [7:0] n1372_o;
  wire [31:0] n1373_o;
  wire n1374_o;
  wire [4:0] n1375_o;
  wire n1376_o;
  wire [11:0] n1377_o;
  wire n1378_o;
  wire [3:0] n1379_o;
  wire [63:0] n1380_o;
  wire [63:0] n1381_o;
  wire n1382_o;
  wire n1383_o;
  wire n1384_o;
  wire [15:0] n1385_o;
  wire [63:0] n1386_o;
  wire n1387_o;
  wire [2:0] n1388_o;
  wire n1389_o;
  wire [6:0] n1390_o;
  wire [63:0] n1391_o;
  wire [4:0] n1392_o;
  wire n1393_o;
  wire n1394_o;
  wire n1395_o;
  wire [11:0] n1396_o;
  wire [63:0] n1397_o;
  wire [15:0] n1398_o;
  wire n1399_o;
  wire n1400_o;
  wire [2:0] n1401_o;
  wire n1402_o;
  wire [6:0] n1403_o;
  wire [63:0] n1404_o;
  wire n1405_o;
  wire [7:0] n1406_o;
  wire [31:0] n1407_o;
  wire [11:0] n1408_o;
  wire [63:0] n1409_o;
  wire [15:0] n1410_o;
  wire [71:0] n1411_o;
  wire [46:0] n1413_o;
  wire [134:0] n1415_o;
  wire [1:0] n1417_o;
  wire [2:0] n1421_o;
  wire [63:0] debug_0_dmi_dout;
  wire debug_0_dmi_ack;
  wire debug_0_core_stop;
  wire debug_0_core_rst;
  wire debug_0_icache_rst;
  wire debug_0_dbg_gpr_req;
  wire [6:0] debug_0_dbg_gpr_addr;
  wire [63:0] debug_0_log_read_data;
  wire [31:0] debug_0_log_write_addr;
  wire debug_0_terminated_out;
  wire [63:0] n1430_o;
  reg n1437_q;
  reg n1439_q;
  reg n1440_q;
  reg n1441_q;
  reg n1442_q;
  reg n1443_q;
  reg n1444_q;
  reg n1445_q;
  reg n1446_q;
  reg n1447_q;
  reg n1448_q;
  wire [255:0] n1449_o;
  assign wishbone_insn_out_adr = n1006_o;
  assign wishbone_insn_out_dat = n1007_o;
  assign wishbone_insn_out_sel = n1008_o;
  assign wishbone_insn_out_cyc = n1009_o;
  assign wishbone_insn_out_stb = n1010_o;
  assign wishbone_insn_out_we = n1011_o;
  assign wishbone_data_out_adr = n1014_o;
  assign wishbone_data_out_dat = n1015_o;
  assign wishbone_data_out_sel = n1016_o;
  assign wishbone_data_out_cyc = n1017_o;
  assign wishbone_data_out_stb = n1018_o;
  assign wishbone_data_out_we = n1019_o;
  assign dmi_dout = debug_0_dmi_dout;
  assign dmi_ack = debug_0_dmi_ack;
  assign terminated_out = debug_0_terminated_out;
  /* soc.vhdl:1096:28  */
  assign n1004_o = {wishbone_insn_in_stall, wishbone_insn_in_ack, wishbone_insn_in_dat};
  /* soc.vhdl:1090:30  */
  assign n1006_o = n1086_o[28:0];
  /* soc.vhdl:1016:30  */
  assign n1007_o = n1086_o[92:29];
  /* soc.vhdl:1010:28  */
  assign n1008_o = n1086_o[100:93];
  /* soc.vhdl:1009:36  */
  assign n1009_o = n1086_o[101];
  /* soc.vhdl:1008:36  */
  assign n1010_o = n1086_o[102];
  /* soc.vhdl:1006:36  */
  assign n1011_o = n1086_o[103];
  /* soc.vhdl:986:33  */
  assign n1012_o = {wishbone_data_in_stall, wishbone_data_in_ack, wishbone_data_in_dat};
  /* soc.vhdl:959:29  */
  assign n1014_o = n1356_o[28:0];
  /* soc.vhdl:958:29  */
  assign n1015_o = n1356_o[92:29];
  /* soc.vhdl:956:29  */
  assign n1016_o = n1356_o[100:93];
  /* soc.vhdl:944:24  */
  assign n1017_o = n1356_o[101];
  /* soc.vhdl:942:23  */
  assign n1018_o = n1356_o[102];
  /* soc.vhdl:930:29  */
  assign n1019_o = n1356_o[103];
  /* soc.vhdl:928:23  */
  assign n1020_o = {wb_snoop_in_we, wb_snoop_in_stb, wb_snoop_in_cyc, wb_snoop_in_sel, wb_snoop_in_dat, wb_snoop_in_adr};
  /* core.vhdl:58:12  */
  assign fetch1_to_icache = n1064_o; // (signal)
  /* core.vhdl:59:12  */
  assign writeback_to_fetch1 = n1415_o; // (signal)
  /* core.vhdl:60:12  */
  assign icache_to_decode1 = n1077_o; // (signal)
  /* core.vhdl:61:12  */
  assign mmu_to_icache = n1324_o; // (signal)
  /* core.vhdl:64:12  */
  assign decode1_to_decode2 = n1112_o; // (signal)
  /* core.vhdl:65:12  */
  assign decode1_to_fetch1 = n1110_o; // (signal)
  /* core.vhdl:66:12  */
  assign decode2_to_execute1 = n1129_o; // (signal)
  /* core.vhdl:69:12  */
  assign register_file_to_decode2 = n1150_o; // (signal)
  /* core.vhdl:70:12  */
  assign decode2_to_register_file = n1134_o; // (signal)
  /* core.vhdl:71:12  */
  assign writeback_to_register_file = n1411_o; // (signal)
  /* core.vhdl:74:12  */
  assign decode2_to_cr_file = decode2_0_c_out_read; // (signal)
  /* core.vhdl:75:12  */
  assign cr_file_to_decode2 = n1160_o; // (signal)
  /* core.vhdl:76:12  */
  assign writeback_to_cr_file = n1413_o; // (signal)
  /* core.vhdl:79:12  */
  assign execute1_to_writeback = n1218_o; // (signal)
  /* core.vhdl:80:12  */
  assign execute1_bypass = n1220_o; // (signal)
  /* core.vhdl:81:12  */
  assign execute1_cr_bypass = n1222_o; // (signal)
  /* core.vhdl:84:12  */
  assign execute1_to_loadstore1 = n1214_o; // (signal)
  /* core.vhdl:85:12  */
  assign loadstore1_to_execute1 = n1282_o; // (signal)
  /* core.vhdl:86:12  */
  assign loadstore1_to_writeback = n1284_o; // (signal)
  /* core.vhdl:87:12  */
  assign loadstore1_to_mmu = n1293_o; // (signal)
  /* core.vhdl:88:12  */
  assign mmu_to_loadstore1 = n1316_o; // (signal)
  /* core.vhdl:91:12  */
  assign loadstore1_to_dcache = n1286_o; // (signal)
  /* core.vhdl:92:12  */
  assign dcache_to_loadstore1 = n1339_o; // (signal)
  /* core.vhdl:93:12  */
  assign mmu_to_dcache = n1318_o; // (signal)
  /* core.vhdl:94:12  */
  assign dcache_to_mmu = n1347_o; // (signal)
  /* core.vhdl:97:12  */
  assign execute1_to_fpu = n1216_o; // (signal)
  /* core.vhdl:98:12  */
  assign fpu_to_execute1 = n1254_o; // (signal)
  /* core.vhdl:99:12  */
  assign fpu_to_writeback = n1256_o; // (signal)
  /* core.vhdl:102:12  */
  assign fetch1_stall_in = n1067_o; // (signal)
  /* core.vhdl:103:12  */
  assign icache_stall_out = icache_0_stall_out; // (signal)
  /* core.vhdl:104:12  */
  assign icache_stall_in = decode1_busy; // (signal)
  /* core.vhdl:105:12  */
  assign decode1_stall_in = decode2_stall_out; // (signal)
  /* core.vhdl:106:12  */
  assign decode1_busy = decode1_0_busy_out; // (signal)
  /* core.vhdl:107:12  */
  assign decode2_busy_in = ex1_busy_out; // (signal)
  /* core.vhdl:108:12  */
  assign decode2_stall_out = decode2_0_stall_out; // (signal)
  /* core.vhdl:109:12  */
  assign ex1_icache_inval = execute1_0_icache_inval; // (signal)
  /* core.vhdl:110:12  */
  assign ex1_busy_out = execute1_0_busy_out; // (signal)
  /* core.vhdl:111:12  */
  assign dcache_stall_out = dcache_0_stall_out; // (signal)
  /* core.vhdl:113:12  */
  assign flush = writeback_0_flush_out; // (signal)
  /* core.vhdl:114:12  */
  assign decode1_flush = decode1_0_flush_out; // (signal)
  /* core.vhdl:115:12  */
  assign fetch1_flush = n1068_o; // (signal)
  /* core.vhdl:117:12  */
  assign complete = n1421_o; // (signal)
  /* core.vhdl:118:12  */
  assign terminate = execute1_0_terminate_out; // (signal)
  /* core.vhdl:119:12  */
  assign core_rst = n1035_o; // (signal)
  /* core.vhdl:121:12  */
  assign do_interrupt = writeback_0_interrupt_out; // (signal)
  /* core.vhdl:124:12  */
  always @*
    rst_fetch1 = n1437_q; // (isignal)
  initial
    rst_fetch1 = 1'b1;
  /* core.vhdl:126:12  */
  always @*
    rst_icache = n1439_q; // (isignal)
  initial
    rst_icache = 1'b1;
  /* core.vhdl:127:12  */
  always @*
    rst_dcache = n1440_q; // (isignal)
  initial
    rst_dcache = 1'b1;
  /* core.vhdl:128:12  */
  always @*
    rst_dec1 = n1441_q; // (isignal)
  initial
    rst_dec1 = 1'b1;
  /* core.vhdl:129:12  */
  always @*
    rst_dec2 = n1442_q; // (isignal)
  initial
    rst_dec2 = 1'b1;
  /* core.vhdl:130:12  */
  always @*
    rst_ex1 = n1443_q; // (isignal)
  initial
    rst_ex1 = 1'b1;
  /* core.vhdl:131:12  */
  always @*
    rst_fpu = n1444_q; // (isignal)
  initial
    rst_fpu = 1'b1;
  /* core.vhdl:132:12  */
  always @*
    rst_ls1 = n1445_q; // (isignal)
  initial
    rst_ls1 = 1'b1;
  /* core.vhdl:133:12  */
  always @*
    rst_wback = n1446_q; // (isignal)
  initial
    rst_wback = 1'b1;
  /* core.vhdl:134:12  */
  always @*
    rst_dbg = n1447_q; // (isignal)
  initial
    rst_dbg = 1'b1;
  /* core.vhdl:135:12  */
  assign alt_reset_d = n1448_q; // (signal)
  /* core.vhdl:137:12  */
  assign sim_cr_dump = register_file_0_sim_dump_done; // (signal)
  /* core.vhdl:140:12  */
  assign dbg_core_stop = debug_0_core_stop; // (signal)
  /* core.vhdl:141:12  */
  assign dbg_core_rst = debug_0_core_rst; // (signal)
  /* core.vhdl:142:12  */
  assign dbg_icache_rst = debug_0_icache_rst; // (signal)
  /* core.vhdl:144:12  */
  assign dbg_gpr_req = debug_0_dbg_gpr_req; // (signal)
  /* core.vhdl:145:12  */
  assign dbg_gpr_ack = register_file_0_dbg_gpr_ack; // (signal)
  /* core.vhdl:146:12  */
  assign dbg_gpr_addr = debug_0_dbg_gpr_addr; // (signal)
  /* core.vhdl:147:12  */
  assign dbg_gpr_data = register_file_0_dbg_gpr_data; // (signal)
  /* core.vhdl:149:12  */
  assign msr = execute1_0_dbg_msr_out; // (signal)
  /* core.vhdl:152:12  */
  assign icache_events = n1097_o; // (signal)
  /* core.vhdl:153:12  */
  assign loadstore_events = n1303_o; // (signal)
  /* core.vhdl:154:12  */
  assign dcache_events = n1361_o; // (signal)
  /* core.vhdl:155:12  */
  assign writeback_events = n1417_o; // (signal)
  /* core.vhdl:158:12  */
  assign dbg_core_is_stopped = decode2_0_stopped_out; // (signal)
  /* core.vhdl:161:12  */
  assign log_data = n1449_o; // (signal)
  /* core.vhdl:162:12  */
  assign log_rd_addr = execute1_0_log_rd_addr; // (signal)
  /* core.vhdl:163:12  */
  assign log_wr_addr = debug_0_log_write_addr; // (signal)
  /* core.vhdl:164:12  */
  assign log_rd_data = debug_0_log_read_data; // (signal)
  /* core.vhdl:189:30  */
  assign n1035_o = dbg_core_rst | rst;
  /* core.vhdl:209:5  */
  fetch1_1e2926114d55612f17be0ce20b92717fa98c0d5f fetch1_0 (
    .clk(clk),
    .rst(rst_fetch1),
    .stall_in(fetch1_stall_in),
    .flush_in(fetch1_flush),
    .inval_btc(n1052_o),
    .stop_in(dbg_core_stop),
    .alt_reset_in(alt_reset_d),
    .w_in_redirect(n1053_o),
    .w_in_virt_mode(n1054_o),
    .w_in_priv_mode(n1055_o),
    .w_in_big_endian(n1056_o),
    .w_in_mode_32bit(n1057_o),
    .w_in_redirect_nia(n1058_o),
    .w_in_br_nia(n1059_o),
    .w_in_br_last(n1060_o),
    .w_in_br_taken(n1061_o),
    .d_in_redirect(n1062_o),
    .d_in_redirect_nia(n1063_o),
    .i_out_req(fetch1_0_i_out_req),
    .i_out_virt_mode(fetch1_0_i_out_virt_mode),
    .i_out_priv_mode(fetch1_0_i_out_priv_mode),
    .i_out_big_endian(fetch1_0_i_out_big_endian),
    .i_out_stop_mark(fetch1_0_i_out_stop_mark),
    .i_out_predicted(fetch1_0_i_out_predicted),
    .i_out_pred_ntaken(fetch1_0_i_out_pred_ntaken),
    .i_out_nia(fetch1_0_i_out_nia),
    .log_out(fetch1_0_log_out));
  /* core.vhdl:221:60  */
  assign n1051_o = mmu_to_icache[1];
  /* core.vhdl:221:43  */
  assign n1052_o = ex1_icache_inval | n1051_o;
  /* soc.vhdl:402:5  */
  assign n1053_o = writeback_to_fetch1[0];
  assign n1054_o = writeback_to_fetch1[1];
  assign n1055_o = writeback_to_fetch1[2];
  assign n1056_o = writeback_to_fetch1[3];
  /* soc.vhdl:285:18  */
  assign n1057_o = writeback_to_fetch1[4];
  assign n1058_o = writeback_to_fetch1[68:5];
  /* soc.vhdl:283:14  */
  assign n1059_o = writeback_to_fetch1[132:69];
  /* soc.vhdl:283:14  */
  assign n1060_o = writeback_to_fetch1[133];
  assign n1061_o = writeback_to_fetch1[134];
  /* soc.vhdl:283:14  */
  assign n1062_o = decode1_to_fetch1[0];
  assign n1063_o = decode1_to_fetch1[64:1];
  assign n1064_o = {fetch1_0_i_out_nia, fetch1_0_i_out_pred_ntaken, fetch1_0_i_out_predicted, fetch1_0_i_out_stop_mark, fetch1_0_i_out_big_endian, fetch1_0_i_out_priv_mode, fetch1_0_i_out_virt_mode, fetch1_0_i_out_req};
  /* core.vhdl:229:41  */
  assign n1067_o = icache_stall_out | decode1_busy;
  /* core.vhdl:230:27  */
  assign n1068_o = flush | decode1_flush;
  /* core.vhdl:232:5  */
  icache_64_8_4_1_4_12_0_5ba93c9db0cff93f52b521d7420e43f6eda2784f icache_0 (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(clk),
    .rst(rst_icache),
    .i_in_req(n1069_o),
    .i_in_virt_mode(n1070_o),
    .i_in_priv_mode(n1071_o),
    .i_in_big_endian(n1072_o),
    .i_in_stop_mark(n1073_o),
    .i_in_predicted(n1074_o),
    .i_in_pred_ntaken(n1075_o),
    .i_in_nia(n1076_o),
    .m_in_tlbld(n1079_o),
    .m_in_tlbie(n1080_o),
    .m_in_doall(n1081_o),
    .m_in_addr(n1082_o),
    .m_in_pte(n1083_o),
    .stall_in(icache_stall_in),
    .flush_in(fetch1_flush),
    .inval_in(n1085_o),
    .wishbone_in_dat(n1088_o),
    .wishbone_in_ack(n1089_o),
    .wishbone_in_stall(n1090_o),
    .wb_snoop_in_adr(n1091_o),
    .wb_snoop_in_dat(n1092_o),
    .wb_snoop_in_sel(n1093_o),
    .wb_snoop_in_cyc(n1094_o),
    .wb_snoop_in_stb(n1095_o),
    .wb_snoop_in_we(n1096_o),
    .i_out_valid(icache_0_i_out_valid),
    .i_out_stop_mark(icache_0_i_out_stop_mark),
    .i_out_fetch_failed(icache_0_i_out_fetch_failed),
    .i_out_nia(icache_0_i_out_nia),
    .i_out_insn(icache_0_i_out_insn),
    .i_out_big_endian(icache_0_i_out_big_endian),
    .i_out_next_predicted(icache_0_i_out_next_predicted),
    .i_out_next_pred_ntaken(icache_0_i_out_next_pred_ntaken),
    .stall_out(icache_0_stall_out),
    .wishbone_out_adr(icache_0_wishbone_out_adr),
    .wishbone_out_dat(icache_0_wishbone_out_dat),
    .wishbone_out_sel(icache_0_wishbone_out_sel),
    .wishbone_out_cyc(icache_0_wishbone_out_cyc),
    .wishbone_out_stb(icache_0_wishbone_out_stb),
    .wishbone_out_we(icache_0_wishbone_out_we),
    .events_icache_miss(icache_0_events_icache_miss),
    .events_itlb_miss_resolved(icache_0_events_itlb_miss_resolved),
    .log_out(icache_0_log_out));
  /* soc.vhdl:267:18  */
  assign n1069_o = fetch1_to_icache[0];
  assign n1070_o = fetch1_to_icache[1];
  /* soc.vhdl:266:14  */
  assign n1071_o = fetch1_to_icache[2];
  /* soc.vhdl:266:14  */
  assign n1072_o = fetch1_to_icache[3];
  assign n1073_o = fetch1_to_icache[4];
  /* soc.vhdl:266:14  */
  assign n1074_o = fetch1_to_icache[5];
  assign n1075_o = fetch1_to_icache[6];
  /* soc.vhdl:324:5  */
  assign n1076_o = fetch1_to_icache[70:7];
  /* soc.vhdl:190:12  */
  assign n1077_o = {icache_0_i_out_next_pred_ntaken, icache_0_i_out_next_predicted, icache_0_i_out_big_endian, icache_0_i_out_insn, icache_0_i_out_nia, icache_0_i_out_fetch_failed, icache_0_i_out_stop_mark, icache_0_i_out_valid};
  assign n1079_o = mmu_to_icache[0];
  assign n1080_o = mmu_to_icache[1];
  assign n1081_o = mmu_to_icache[2];
  assign n1082_o = mmu_to_icache[66:3];
  assign n1083_o = mmu_to_icache[130:67];
  /* core.vhdl:248:40  */
  assign n1085_o = dbg_icache_rst | ex1_icache_inval;
  assign n1086_o = {icache_0_wishbone_out_we, icache_0_wishbone_out_stb, icache_0_wishbone_out_cyc, icache_0_wishbone_out_sel, icache_0_wishbone_out_dat, icache_0_wishbone_out_adr};
  assign n1088_o = n1004_o[63:0];
  assign n1089_o = n1004_o[64];
  assign n1090_o = n1004_o[65];
  assign n1091_o = n1020_o[28:0];
  assign n1092_o = n1020_o[92:29];
  assign n1093_o = n1020_o[100:93];
  assign n1094_o = n1020_o[101];
  assign n1095_o = n1020_o[102];
  assign n1096_o = n1020_o[103];
  assign n1097_o = {icache_0_events_itlb_miss_resolved, icache_0_events_icache_miss};
  /* core.vhdl:260:5  */
  decode1_0_bf8b4530d8d246dd74ac53a13471bba17941dff7 decode1_0 (
    .clk(clk),
    .rst(rst_dec1),
    .stall_in(decode1_stall_in),
    .flush_in(flush),
    .f_in_valid(n1102_o),
    .f_in_stop_mark(n1103_o),
    .f_in_fetch_failed(n1104_o),
    .f_in_nia(n1105_o),
    .f_in_insn(n1106_o),
    .f_in_big_endian(n1107_o),
    .f_in_next_predicted(n1108_o),
    .f_in_next_pred_ntaken(n1109_o),
    .busy_out(decode1_0_busy_out),
    .flush_out(decode1_0_flush_out),
    .f_out_redirect(decode1_0_f_out_redirect),
    .f_out_redirect_nia(decode1_0_f_out_redirect_nia),
    .d_out_valid(decode1_0_d_out_valid),
    .d_out_stop_mark(decode1_0_d_out_stop_mark),
    .d_out_nia(decode1_0_d_out_nia),
    .d_out_insn(decode1_0_d_out_insn),
    .d_out_ispr1(decode1_0_d_out_ispr1),
    .d_out_ispr2(decode1_0_d_out_ispr2),
    .d_out_ispro(decode1_0_d_out_ispro),
    .d_out_decode(decode1_0_d_out_decode),
    .d_out_br_pred(decode1_0_d_out_br_pred),
    .d_out_big_endian(decode1_0_d_out_big_endian),
    .log_out(decode1_0_log_out));
  assign n1102_o = icache_to_decode1[0];
  assign n1103_o = icache_to_decode1[1];
  assign n1104_o = icache_to_decode1[2];
  assign n1105_o = icache_to_decode1[66:3];
  assign n1106_o = icache_to_decode1[98:67];
  assign n1107_o = icache_to_decode1[99];
  assign n1108_o = icache_to_decode1[100];
  assign n1109_o = icache_to_decode1[101];
  assign n1110_o = {decode1_0_f_out_redirect_nia, decode1_0_f_out_redirect};
  assign n1112_o = {decode1_0_d_out_big_endian, decode1_0_d_out_br_pred, decode1_0_d_out_decode, decode1_0_d_out_ispro, decode1_0_d_out_ispr2, decode1_0_d_out_ispr1, decode1_0_d_out_insn, decode1_0_d_out_nia, decode1_0_d_out_stop_mark, decode1_0_d_out_valid};
  /* core.vhdl:280:5  */
  decode2_0_9159cb8bcee7fcb95582f140960cdae72788d326 decode2_0 (
    .clk(clk),
    .rst(rst_dec2),
    .complete_in_tag(n1115_o),
    .complete_in_valid(n1116_o),
    .busy_in(decode2_busy_in),
    .flush_in(flush),
    .d_in_valid(n1119_o),
    .d_in_stop_mark(n1120_o),
    .d_in_nia(n1121_o),
    .d_in_insn(n1122_o),
    .d_in_ispr1(n1123_o),
    .d_in_ispr2(n1124_o),
    .d_in_ispro(n1125_o),
    .d_in_decode(n1126_o),
    .d_in_br_pred(n1127_o),
    .d_in_big_endian(n1128_o),
    .r_in_read1_data(n1131_o),
    .r_in_read2_data(n1132_o),
    .r_in_read3_data(n1133_o),
    .c_in_read_cr_data(n1136_o),
    .c_in_read_xerc_data(n1137_o),
    .execute_bypass_tag(n1139_o),
    .execute_bypass_data(n1140_o),
    .execute_cr_bypass_tag(n1141_o),
    .execute_cr_bypass_data(n1142_o),
    .stall_out(decode2_0_stall_out),
    .stopped_out(decode2_0_stopped_out),
    .e_out_valid(decode2_0_e_out_valid),
    .e_out_unit(decode2_0_e_out_unit),
    .e_out_fac(decode2_0_e_out_fac),
    .e_out_insn_type(decode2_0_e_out_insn_type),
    .e_out_nia(decode2_0_e_out_nia),
    .e_out_instr_tag(decode2_0_e_out_instr_tag),
    .e_out_write_reg(decode2_0_e_out_write_reg),
    .e_out_write_reg_enable(decode2_0_e_out_write_reg_enable),
    .e_out_read_reg1(decode2_0_e_out_read_reg1),
    .e_out_read_reg2(decode2_0_e_out_read_reg2),
    .e_out_read_data1(decode2_0_e_out_read_data1),
    .e_out_read_data2(decode2_0_e_out_read_data2),
    .e_out_read_data3(decode2_0_e_out_read_data3),
    .e_out_cr(decode2_0_e_out_cr),
    .e_out_xerc(decode2_0_e_out_xerc),
    .e_out_lr(decode2_0_e_out_lr),
    .e_out_br_abs(decode2_0_e_out_br_abs),
    .e_out_rc(decode2_0_e_out_rc),
    .e_out_oe(decode2_0_e_out_oe),
    .e_out_invert_a(decode2_0_e_out_invert_a),
    .e_out_addm1(decode2_0_e_out_addm1),
    .e_out_invert_out(decode2_0_e_out_invert_out),
    .e_out_input_carry(decode2_0_e_out_input_carry),
    .e_out_output_carry(decode2_0_e_out_output_carry),
    .e_out_input_cr(decode2_0_e_out_input_cr),
    .e_out_output_cr(decode2_0_e_out_output_cr),
    .e_out_output_xer(decode2_0_e_out_output_xer),
    .e_out_is_32bit(decode2_0_e_out_is_32bit),
    .e_out_is_signed(decode2_0_e_out_is_signed),
    .e_out_insn(decode2_0_e_out_insn),
    .e_out_data_len(decode2_0_e_out_data_len),
    .e_out_byte_reverse(decode2_0_e_out_byte_reverse),
    .e_out_sign_extend(decode2_0_e_out_sign_extend),
    .e_out_update(decode2_0_e_out_update),
    .e_out_reserve(decode2_0_e_out_reserve),
    .e_out_br_pred(decode2_0_e_out_br_pred),
    .e_out_result_sel(decode2_0_e_out_result_sel),
    .e_out_sub_select(decode2_0_e_out_sub_select),
    .e_out_repeat(decode2_0_e_out_repeat),
    .e_out_second(decode2_0_e_out_second),
    .r_out_read1_enable(decode2_0_r_out_read1_enable),
    .r_out_read1_reg(decode2_0_r_out_read1_reg),
    .r_out_read2_enable(decode2_0_r_out_read2_enable),
    .r_out_read2_reg(decode2_0_r_out_read2_reg),
    .r_out_read3_enable(decode2_0_r_out_read3_enable),
    .r_out_read3_reg(decode2_0_r_out_read3_reg),
    .c_out_read(decode2_0_c_out_read),
    .log_out(decode2_0_log_out));
  assign n1115_o = complete[1:0];
  assign n1116_o = complete[2];
  assign n1119_o = decode1_to_decode2[0];
  assign n1120_o = decode1_to_decode2[1];
  assign n1121_o = decode1_to_decode2[65:2];
  assign n1122_o = decode1_to_decode2[97:66];
  assign n1123_o = decode1_to_decode2[104:98];
  assign n1124_o = decode1_to_decode2[111:105];
  assign n1125_o = decode1_to_decode2[118:112];
  assign n1126_o = decode1_to_decode2[162:119];
  assign n1127_o = decode1_to_decode2[163];
  assign n1128_o = decode1_to_decode2[164];
  assign n1129_o = {decode2_0_e_out_second, decode2_0_e_out_repeat, decode2_0_e_out_sub_select, decode2_0_e_out_result_sel, decode2_0_e_out_br_pred, decode2_0_e_out_reserve, decode2_0_e_out_update, decode2_0_e_out_sign_extend, decode2_0_e_out_byte_reverse, decode2_0_e_out_data_len, decode2_0_e_out_insn, decode2_0_e_out_is_signed, decode2_0_e_out_is_32bit, decode2_0_e_out_output_xer, decode2_0_e_out_output_cr, decode2_0_e_out_input_cr, decode2_0_e_out_output_carry, decode2_0_e_out_input_carry, decode2_0_e_out_invert_out, decode2_0_e_out_addm1, decode2_0_e_out_invert_a, decode2_0_e_out_oe, decode2_0_e_out_rc, decode2_0_e_out_br_abs, decode2_0_e_out_lr, decode2_0_e_out_xerc, decode2_0_e_out_cr, decode2_0_e_out_read_data3, decode2_0_e_out_read_data2, decode2_0_e_out_read_data1, decode2_0_e_out_read_reg2, decode2_0_e_out_read_reg1, decode2_0_e_out_write_reg_enable, decode2_0_e_out_write_reg, decode2_0_e_out_instr_tag, decode2_0_e_out_nia, decode2_0_e_out_insn_type, decode2_0_e_out_fac, decode2_0_e_out_unit, decode2_0_e_out_valid};
  assign n1131_o = register_file_to_decode2[63:0];
  assign n1132_o = register_file_to_decode2[127:64];
  assign n1133_o = register_file_to_decode2[191:128];
  assign n1134_o = {decode2_0_r_out_read3_reg, decode2_0_r_out_read3_enable, decode2_0_r_out_read2_reg, decode2_0_r_out_read2_enable, decode2_0_r_out_read1_reg, decode2_0_r_out_read1_enable};
  assign n1136_o = cr_file_to_decode2[31:0];
  assign n1137_o = cr_file_to_decode2[36:32];
  assign n1139_o = execute1_bypass[2:0];
  assign n1140_o = execute1_bypass[66:3];
  assign n1141_o = execute1_cr_bypass[2:0];
  assign n1142_o = execute1_cr_bypass[34:3];
  /* core.vhdl:306:5  */
  register_file_0_3f29546453678b855931c174a97d6c0894b8f546 register_file_0 (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(clk),
    .d_in_read1_enable(n1144_o),
    .d_in_read1_reg(n1145_o),
    .d_in_read2_enable(n1146_o),
    .d_in_read2_reg(n1147_o),
    .d_in_read3_enable(n1148_o),
    .d_in_read3_reg(n1149_o),
    .w_in_write_reg(n1152_o),
    .w_in_write_data(n1153_o),
    .w_in_write_enable(n1154_o),
    .dbg_gpr_req(dbg_gpr_req),
    .dbg_gpr_addr(dbg_gpr_addr),
    .sim_dump(terminate),
    .d_out_read1_data(register_file_0_d_out_read1_data),
    .d_out_read2_data(register_file_0_d_out_read2_data),
    .d_out_read3_data(register_file_0_d_out_read3_data),
    .dbg_gpr_ack(register_file_0_dbg_gpr_ack),
    .dbg_gpr_data(register_file_0_dbg_gpr_data),
    .sim_dump_done(register_file_0_sim_dump_done),
    .log_out(register_file_0_log_out));
  assign n1144_o = decode2_to_register_file[0];
  assign n1145_o = decode2_to_register_file[7:1];
  assign n1146_o = decode2_to_register_file[8];
  assign n1147_o = decode2_to_register_file[15:9];
  assign n1148_o = decode2_to_register_file[16];
  assign n1149_o = decode2_to_register_file[23:17];
  assign n1150_o = {register_file_0_d_out_read3_data, register_file_0_d_out_read2_data, register_file_0_d_out_read1_data};
  assign n1152_o = writeback_to_register_file[6:0];
  assign n1153_o = writeback_to_register_file[70:7];
  assign n1154_o = writeback_to_register_file[71];
  /* core.vhdl:326:5  */
  cr_file_0_5ba93c9db0cff93f52b521d7420e43f6eda2784f cr_file_0 (
    .clk(clk),
    .d_in_read(n1159_o),
    .w_in_write_cr_enable(n1162_o),
    .w_in_write_cr_mask(n1163_o),
    .w_in_write_cr_data(n1164_o),
    .w_in_write_xerc_enable(n1165_o),
    .w_in_write_xerc_data(n1166_o),
    .sim_dump(sim_cr_dump),
    .d_out_read_cr_data(cr_file_0_d_out_read_cr_data),
    .d_out_read_xerc_data(cr_file_0_d_out_read_xerc_data),
    .log_out(cr_file_0_log_out));
  assign n1159_o = decode2_to_cr_file;
  assign n1160_o = {cr_file_0_d_out_read_xerc_data, cr_file_0_d_out_read_cr_data};
  assign n1162_o = writeback_to_cr_file[0];
  assign n1163_o = writeback_to_cr_file[8:1];
  assign n1164_o = writeback_to_cr_file[40:9];
  assign n1165_o = writeback_to_cr_file[41];
  assign n1166_o = writeback_to_cr_file[46:42];
  /* core.vhdl:340:5  */
  execute1_0_47ec8d98366433dc002e7721c9e37d5067547937 execute1_0 (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(clk),
    .rst(rst_ex1),
    .flush_in(flush),
    .e_in_valid(n1169_o),
    .e_in_unit(n1170_o),
    .e_in_fac(n1171_o),
    .e_in_insn_type(n1172_o),
    .e_in_nia(n1173_o),
    .e_in_instr_tag(n1174_o),
    .e_in_write_reg(n1175_o),
    .e_in_write_reg_enable(n1176_o),
    .e_in_read_reg1(n1177_o),
    .e_in_read_reg2(n1178_o),
    .e_in_read_data1(n1179_o),
    .e_in_read_data2(n1180_o),
    .e_in_read_data3(n1181_o),
    .e_in_cr(n1182_o),
    .e_in_xerc(n1183_o),
    .e_in_lr(n1184_o),
    .e_in_br_abs(n1185_o),
    .e_in_rc(n1186_o),
    .e_in_oe(n1187_o),
    .e_in_invert_a(n1188_o),
    .e_in_addm1(n1189_o),
    .e_in_invert_out(n1190_o),
    .e_in_input_carry(n1191_o),
    .e_in_output_carry(n1192_o),
    .e_in_input_cr(n1193_o),
    .e_in_output_cr(n1194_o),
    .e_in_output_xer(n1195_o),
    .e_in_is_32bit(n1196_o),
    .e_in_is_signed(n1197_o),
    .e_in_insn(n1198_o),
    .e_in_data_len(n1199_o),
    .e_in_byte_reverse(n1200_o),
    .e_in_sign_extend(n1201_o),
    .e_in_update(n1202_o),
    .e_in_reserve(n1203_o),
    .e_in_br_pred(n1204_o),
    .e_in_result_sel(n1205_o),
    .e_in_sub_select(n1206_o),
    .e_in_repeat(n1207_o),
    .e_in_second(n1208_o),
    .l_in_busy(n1209_o),
    .l_in_in_progress(n1210_o),
    .l_in_interrupt(n1211_o),
    .fp_in_busy(n1212_o),
    .fp_in_exception(n1213_o),
    .ext_irq_in(ext_irq),
    .interrupt_in(do_interrupt),
    .wb_events_instr_complete(n1227_o),
    .wb_events_fp_complete(n1228_o),
    .ls_events_load_complete(n1229_o),
    .ls_events_store_complete(n1230_o),
    .ls_events_itlb_miss(n1231_o),
    .dc_events_load_miss(n1232_o),
    .dc_events_store_miss(n1233_o),
    .dc_events_dcache_refill(n1234_o),
    .dc_events_dtlb_miss(n1235_o),
    .dc_events_dtlb_miss_resolved(n1236_o),
    .ic_events_icache_miss(n1237_o),
    .ic_events_itlb_miss_resolved(n1238_o),
    .log_rd_data(log_rd_data),
    .log_wr_addr(log_wr_addr),
    .busy_out(execute1_0_busy_out),
    .l_out_valid(execute1_0_l_out_valid),
    .l_out_op(execute1_0_l_out_op),
    .l_out_nia(execute1_0_l_out_nia),
    .l_out_insn(execute1_0_l_out_insn),
    .l_out_instr_tag(execute1_0_l_out_instr_tag),
    .l_out_addr1(execute1_0_l_out_addr1),
    .l_out_addr2(execute1_0_l_out_addr2),
    .l_out_data(execute1_0_l_out_data),
    .l_out_write_reg(execute1_0_l_out_write_reg),
    .l_out_length(execute1_0_l_out_length),
    .l_out_ci(execute1_0_l_out_ci),
    .l_out_byte_reverse(execute1_0_l_out_byte_reverse),
    .l_out_sign_extend(execute1_0_l_out_sign_extend),
    .l_out_update(execute1_0_l_out_update),
    .l_out_xerc(execute1_0_l_out_xerc),
    .l_out_reserve(execute1_0_l_out_reserve),
    .l_out_rc(execute1_0_l_out_rc),
    .l_out_virt_mode(execute1_0_l_out_virt_mode),
    .l_out_priv_mode(execute1_0_l_out_priv_mode),
    .l_out_mode_32bit(execute1_0_l_out_mode_32bit),
    .l_out_is_32bit(execute1_0_l_out_is_32bit),
    .l_out_repeat(execute1_0_l_out_repeat),
    .l_out_second(execute1_0_l_out_second),
    .l_out_msr(execute1_0_l_out_msr),
    .fp_out_valid(execute1_0_fp_out_valid),
    .fp_out_op(execute1_0_fp_out_op),
    .fp_out_nia(execute1_0_fp_out_nia),
    .fp_out_itag(execute1_0_fp_out_itag),
    .fp_out_insn(execute1_0_fp_out_insn),
    .fp_out_single(execute1_0_fp_out_single),
    .fp_out_fe_mode(execute1_0_fp_out_fe_mode),
    .fp_out_fra(execute1_0_fp_out_fra),
    .fp_out_frb(execute1_0_fp_out_frb),
    .fp_out_frc(execute1_0_fp_out_frc),
    .fp_out_frt(execute1_0_fp_out_frt),
    .fp_out_rc(execute1_0_fp_out_rc),
    .fp_out_out_cr(execute1_0_fp_out_out_cr),
    .e_out_valid(execute1_0_e_out_valid),
    .e_out_instr_tag(execute1_0_e_out_instr_tag),
    .e_out_rc(execute1_0_e_out_rc),
    .e_out_mode_32bit(execute1_0_e_out_mode_32bit),
    .e_out_write_enable(execute1_0_e_out_write_enable),
    .e_out_write_reg(execute1_0_e_out_write_reg),
    .e_out_write_data(execute1_0_e_out_write_data),
    .e_out_write_cr_enable(execute1_0_e_out_write_cr_enable),
    .e_out_write_cr_mask(execute1_0_e_out_write_cr_mask),
    .e_out_write_cr_data(execute1_0_e_out_write_cr_data),
    .e_out_write_xerc_enable(execute1_0_e_out_write_xerc_enable),
    .e_out_xerc(execute1_0_e_out_xerc),
    .e_out_interrupt(execute1_0_e_out_interrupt),
    .e_out_intr_vec(execute1_0_e_out_intr_vec),
    .e_out_redirect(execute1_0_e_out_redirect),
    .e_out_redir_mode(execute1_0_e_out_redir_mode),
    .e_out_last_nia(execute1_0_e_out_last_nia),
    .e_out_br_offset(execute1_0_e_out_br_offset),
    .e_out_br_last(execute1_0_e_out_br_last),
    .e_out_br_taken(execute1_0_e_out_br_taken),
    .e_out_abs_br(execute1_0_e_out_abs_br),
    .e_out_srr1(execute1_0_e_out_srr1),
    .e_out_msr(execute1_0_e_out_msr),
    .bypass_data_tag(execute1_0_bypass_data_tag),
    .bypass_data_data(execute1_0_bypass_data_data),
    .bypass_cr_data_tag(execute1_0_bypass_cr_data_tag),
    .bypass_cr_data_data(execute1_0_bypass_cr_data_data),
    .dbg_msr_out(execute1_0_dbg_msr_out),
    .icache_inval(execute1_0_icache_inval),
    .terminate_out(execute1_0_terminate_out),
    .log_out(execute1_0_log_out),
    .log_rd_addr(execute1_0_log_rd_addr));
  assign n1169_o = decode2_to_execute1[0];
  assign n1170_o = decode2_to_execute1[2:1];
  assign n1171_o = decode2_to_execute1[3];
  assign n1172_o = decode2_to_execute1[9:4];
  assign n1173_o = decode2_to_execute1[73:10];
  assign n1174_o = decode2_to_execute1[76:74];
  assign n1175_o = decode2_to_execute1[83:77];
  assign n1176_o = decode2_to_execute1[84];
  assign n1177_o = decode2_to_execute1[91:85];
  assign n1178_o = decode2_to_execute1[98:92];
  assign n1179_o = decode2_to_execute1[162:99];
  assign n1180_o = decode2_to_execute1[226:163];
  assign n1181_o = decode2_to_execute1[290:227];
  assign n1182_o = decode2_to_execute1[322:291];
  assign n1183_o = decode2_to_execute1[327:323];
  assign n1184_o = decode2_to_execute1[328];
  assign n1185_o = decode2_to_execute1[329];
  assign n1186_o = decode2_to_execute1[330];
  assign n1187_o = decode2_to_execute1[331];
  assign n1188_o = decode2_to_execute1[332];
  assign n1189_o = decode2_to_execute1[333];
  assign n1190_o = decode2_to_execute1[334];
  assign n1191_o = decode2_to_execute1[336:335];
  assign n1192_o = decode2_to_execute1[337];
  assign n1193_o = decode2_to_execute1[338];
  assign n1194_o = decode2_to_execute1[339];
  assign n1195_o = decode2_to_execute1[340];
  assign n1196_o = decode2_to_execute1[341];
  assign n1197_o = decode2_to_execute1[342];
  assign n1198_o = decode2_to_execute1[374:343];
  assign n1199_o = decode2_to_execute1[378:375];
  assign n1200_o = decode2_to_execute1[379];
  assign n1201_o = decode2_to_execute1[380];
  assign n1202_o = decode2_to_execute1[381];
  assign n1203_o = decode2_to_execute1[382];
  assign n1204_o = decode2_to_execute1[383];
  assign n1205_o = decode2_to_execute1[386:384];
  assign n1206_o = decode2_to_execute1[389:387];
  assign n1207_o = decode2_to_execute1[390];
  assign n1208_o = decode2_to_execute1[391];
  assign n1209_o = loadstore1_to_execute1[0];
  assign n1210_o = loadstore1_to_execute1[1];
  assign n1211_o = loadstore1_to_execute1[2];
  assign n1212_o = fpu_to_execute1[0];
  assign n1213_o = fpu_to_execute1[1];
  assign n1214_o = {execute1_0_l_out_msr, execute1_0_l_out_second, execute1_0_l_out_repeat, execute1_0_l_out_is_32bit, execute1_0_l_out_mode_32bit, execute1_0_l_out_priv_mode, execute1_0_l_out_virt_mode, execute1_0_l_out_rc, execute1_0_l_out_reserve, execute1_0_l_out_xerc, execute1_0_l_out_update, execute1_0_l_out_sign_extend, execute1_0_l_out_byte_reverse, execute1_0_l_out_ci, execute1_0_l_out_length, execute1_0_l_out_write_reg, execute1_0_l_out_data, execute1_0_l_out_addr2, execute1_0_l_out_addr1, execute1_0_l_out_instr_tag, execute1_0_l_out_insn, execute1_0_l_out_nia, execute1_0_l_out_op, execute1_0_l_out_valid};
  assign n1216_o = {execute1_0_fp_out_out_cr, execute1_0_fp_out_rc, execute1_0_fp_out_frt, execute1_0_fp_out_frc, execute1_0_fp_out_frb, execute1_0_fp_out_fra, execute1_0_fp_out_fe_mode, execute1_0_fp_out_single, execute1_0_fp_out_insn, execute1_0_fp_out_itag, execute1_0_fp_out_nia, execute1_0_fp_out_op, execute1_0_fp_out_valid};
  assign n1218_o = {execute1_0_e_out_msr, execute1_0_e_out_srr1, execute1_0_e_out_abs_br, execute1_0_e_out_br_taken, execute1_0_e_out_br_last, execute1_0_e_out_br_offset, execute1_0_e_out_last_nia, execute1_0_e_out_redir_mode, execute1_0_e_out_redirect, execute1_0_e_out_intr_vec, execute1_0_e_out_interrupt, execute1_0_e_out_xerc, execute1_0_e_out_write_xerc_enable, execute1_0_e_out_write_cr_data, execute1_0_e_out_write_cr_mask, execute1_0_e_out_write_cr_enable, execute1_0_e_out_write_data, execute1_0_e_out_write_reg, execute1_0_e_out_write_enable, execute1_0_e_out_mode_32bit, execute1_0_e_out_rc, execute1_0_e_out_instr_tag, execute1_0_e_out_valid};
  assign n1220_o = {execute1_0_bypass_data_data, execute1_0_bypass_data_tag};
  assign n1222_o = {execute1_0_bypass_cr_data_data, execute1_0_bypass_cr_data_tag};
  assign n1227_o = writeback_events[0];
  assign n1228_o = writeback_events[1];
  assign n1229_o = loadstore_events[0];
  assign n1230_o = loadstore_events[1];
  assign n1231_o = loadstore_events[2];
  assign n1232_o = dcache_events[0];
  assign n1233_o = dcache_events[1];
  assign n1234_o = dcache_events[2];
  assign n1235_o = dcache_events[3];
  assign n1236_o = dcache_events[4];
  assign n1237_o = icache_events[0];
  assign n1238_o = icache_events[1];
  /* core.vhdl:377:9  */
  fpu with_fpu_fpu_0 (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(clk),
    .rst(rst_fpu),
    .e_in_valid(n1241_o),
    .e_in_op(n1242_o),
    .e_in_nia(n1243_o),
    .e_in_itag(n1244_o),
    .e_in_insn(n1245_o),
    .e_in_single(n1246_o),
    .e_in_fe_mode(n1247_o),
    .e_in_fra(n1248_o),
    .e_in_frb(n1249_o),
    .e_in_frc(n1250_o),
    .e_in_frt(n1251_o),
    .e_in_rc(n1252_o),
    .e_in_out_cr(n1253_o),
    .e_out_busy(with_fpu_fpu_0_e_out_busy),
    .e_out_exception(with_fpu_fpu_0_e_out_exception),
    .w_out_valid(with_fpu_fpu_0_w_out_valid),
    .w_out_interrupt(with_fpu_fpu_0_w_out_interrupt),
    .w_out_instr_tag(with_fpu_fpu_0_w_out_instr_tag),
    .w_out_write_enable(with_fpu_fpu_0_w_out_write_enable),
    .w_out_write_reg(with_fpu_fpu_0_w_out_write_reg),
    .w_out_write_data(with_fpu_fpu_0_w_out_write_data),
    .w_out_write_cr_enable(with_fpu_fpu_0_w_out_write_cr_enable),
    .w_out_write_cr_mask(with_fpu_fpu_0_w_out_write_cr_mask),
    .w_out_write_cr_data(with_fpu_fpu_0_w_out_write_cr_data),
    .w_out_intr_vec(with_fpu_fpu_0_w_out_intr_vec),
    .w_out_srr0(with_fpu_fpu_0_w_out_srr0),
    .w_out_srr1(with_fpu_fpu_0_w_out_srr1));
  assign n1241_o = execute1_to_fpu[0];
  assign n1242_o = execute1_to_fpu[6:1];
  assign n1243_o = execute1_to_fpu[70:7];
  assign n1244_o = execute1_to_fpu[73:71];
  assign n1245_o = execute1_to_fpu[105:74];
  assign n1246_o = execute1_to_fpu[106];
  assign n1247_o = execute1_to_fpu[108:107];
  assign n1248_o = execute1_to_fpu[172:109];
  assign n1249_o = execute1_to_fpu[236:173];
  assign n1250_o = execute1_to_fpu[300:237];
  assign n1251_o = execute1_to_fpu[307:301];
  assign n1252_o = execute1_to_fpu[308];
  assign n1253_o = execute1_to_fpu[309];
  assign n1254_o = {with_fpu_fpu_0_e_out_exception, with_fpu_fpu_0_e_out_busy};
  assign n1256_o = {with_fpu_fpu_0_w_out_srr1, with_fpu_fpu_0_w_out_srr0, with_fpu_fpu_0_w_out_intr_vec, with_fpu_fpu_0_w_out_write_cr_data, with_fpu_fpu_0_w_out_write_cr_mask, with_fpu_fpu_0_w_out_write_cr_enable, with_fpu_fpu_0_w_out_write_data, with_fpu_fpu_0_w_out_write_reg, with_fpu_fpu_0_w_out_write_enable, with_fpu_fpu_0_w_out_instr_tag, with_fpu_fpu_0_w_out_interrupt, with_fpu_fpu_0_w_out_valid};
  /* core.vhdl:393:5  */
  loadstore1_0_bf8b4530d8d246dd74ac53a13471bba17941dff7 loadstore1_0 (
    .clk(clk),
    .rst(rst_ls1),
    .l_in_valid(n1258_o),
    .l_in_op(n1259_o),
    .l_in_nia(n1260_o),
    .l_in_insn(n1261_o),
    .l_in_instr_tag(n1262_o),
    .l_in_addr1(n1263_o),
    .l_in_addr2(n1264_o),
    .l_in_data(n1265_o),
    .l_in_write_reg(n1266_o),
    .l_in_length(n1267_o),
    .l_in_ci(n1268_o),
    .l_in_byte_reverse(n1269_o),
    .l_in_sign_extend(n1270_o),
    .l_in_update(n1271_o),
    .l_in_xerc(n1272_o),
    .l_in_reserve(n1273_o),
    .l_in_rc(n1274_o),
    .l_in_virt_mode(n1275_o),
    .l_in_priv_mode(n1276_o),
    .l_in_mode_32bit(n1277_o),
    .l_in_is_32bit(n1278_o),
    .l_in_repeat(n1279_o),
    .l_in_second(n1280_o),
    .l_in_msr(n1281_o),
    .d_in_valid(n1288_o),
    .d_in_data(n1289_o),
    .d_in_store_done(n1290_o),
    .d_in_error(n1291_o),
    .d_in_cache_paradox(n1292_o),
    .m_in_done(n1295_o),
    .m_in_err(n1296_o),
    .m_in_invalid(n1297_o),
    .m_in_badtree(n1298_o),
    .m_in_segerr(n1299_o),
    .m_in_perm_error(n1300_o),
    .m_in_rc_error(n1301_o),
    .m_in_sprval(n1302_o),
    .dc_stall(dcache_stall_out),
    .e_out_busy(loadstore1_0_e_out_busy),
    .e_out_in_progress(loadstore1_0_e_out_in_progress),
    .e_out_interrupt(loadstore1_0_e_out_interrupt),
    .l_out_valid(loadstore1_0_l_out_valid),
    .l_out_instr_tag(loadstore1_0_l_out_instr_tag),
    .l_out_write_enable(loadstore1_0_l_out_write_enable),
    .l_out_write_reg(loadstore1_0_l_out_write_reg),
    .l_out_write_data(loadstore1_0_l_out_write_data),
    .l_out_xerc(loadstore1_0_l_out_xerc),
    .l_out_rc(loadstore1_0_l_out_rc),
    .l_out_store_done(loadstore1_0_l_out_store_done),
    .l_out_interrupt(loadstore1_0_l_out_interrupt),
    .l_out_intr_vec(loadstore1_0_l_out_intr_vec),
    .l_out_srr0(loadstore1_0_l_out_srr0),
    .l_out_srr1(loadstore1_0_l_out_srr1),
    .d_out_valid(loadstore1_0_d_out_valid),
    .d_out_hold(loadstore1_0_d_out_hold),
    .d_out_load(loadstore1_0_d_out_load),
    .d_out_dcbz(loadstore1_0_d_out_dcbz),
    .d_out_nc(loadstore1_0_d_out_nc),
    .d_out_reserve(loadstore1_0_d_out_reserve),
    .d_out_atomic(loadstore1_0_d_out_atomic),
    .d_out_atomic_last(loadstore1_0_d_out_atomic_last),
    .d_out_virt_mode(loadstore1_0_d_out_virt_mode),
    .d_out_priv_mode(loadstore1_0_d_out_priv_mode),
    .d_out_addr(loadstore1_0_d_out_addr),
    .d_out_data(loadstore1_0_d_out_data),
    .d_out_byte_sel(loadstore1_0_d_out_byte_sel),
    .m_out_valid(loadstore1_0_m_out_valid),
    .m_out_tlbie(loadstore1_0_m_out_tlbie),
    .m_out_slbia(loadstore1_0_m_out_slbia),
    .m_out_mtspr(loadstore1_0_m_out_mtspr),
    .m_out_iside(loadstore1_0_m_out_iside),
    .m_out_load(loadstore1_0_m_out_load),
    .m_out_priv(loadstore1_0_m_out_priv),
    .m_out_sprn(loadstore1_0_m_out_sprn),
    .m_out_addr(loadstore1_0_m_out_addr),
    .m_out_rs(loadstore1_0_m_out_rs),
    .events_load_complete(loadstore1_0_events_load_complete),
    .events_store_complete(loadstore1_0_events_store_complete),
    .events_itlb_miss(loadstore1_0_events_itlb_miss),
    .log_out(loadstore1_0_log_out));
  assign n1258_o = execute1_to_loadstore1[0];
  assign n1259_o = execute1_to_loadstore1[6:1];
  assign n1260_o = execute1_to_loadstore1[70:7];
  assign n1261_o = execute1_to_loadstore1[102:71];
  assign n1262_o = execute1_to_loadstore1[105:103];
  assign n1263_o = execute1_to_loadstore1[169:106];
  assign n1264_o = execute1_to_loadstore1[233:170];
  assign n1265_o = execute1_to_loadstore1[297:234];
  assign n1266_o = execute1_to_loadstore1[304:298];
  assign n1267_o = execute1_to_loadstore1[308:305];
  assign n1268_o = execute1_to_loadstore1[309];
  assign n1269_o = execute1_to_loadstore1[310];
  assign n1270_o = execute1_to_loadstore1[311];
  assign n1271_o = execute1_to_loadstore1[312];
  assign n1272_o = execute1_to_loadstore1[317:313];
  assign n1273_o = execute1_to_loadstore1[318];
  assign n1274_o = execute1_to_loadstore1[319];
  assign n1275_o = execute1_to_loadstore1[320];
  assign n1276_o = execute1_to_loadstore1[321];
  assign n1277_o = execute1_to_loadstore1[322];
  assign n1278_o = execute1_to_loadstore1[323];
  assign n1279_o = execute1_to_loadstore1[324];
  assign n1280_o = execute1_to_loadstore1[325];
  assign n1281_o = execute1_to_loadstore1[389:326];
  assign n1282_o = {loadstore1_0_e_out_interrupt, loadstore1_0_e_out_in_progress, loadstore1_0_e_out_busy};
  assign n1284_o = {loadstore1_0_l_out_srr1, loadstore1_0_l_out_srr0, loadstore1_0_l_out_intr_vec, loadstore1_0_l_out_interrupt, loadstore1_0_l_out_store_done, loadstore1_0_l_out_rc, loadstore1_0_l_out_xerc, loadstore1_0_l_out_write_data, loadstore1_0_l_out_write_reg, loadstore1_0_l_out_write_enable, loadstore1_0_l_out_instr_tag, loadstore1_0_l_out_valid};
  assign n1286_o = {loadstore1_0_d_out_byte_sel, loadstore1_0_d_out_data, loadstore1_0_d_out_addr, loadstore1_0_d_out_priv_mode, loadstore1_0_d_out_virt_mode, loadstore1_0_d_out_atomic_last, loadstore1_0_d_out_atomic, loadstore1_0_d_out_reserve, loadstore1_0_d_out_nc, loadstore1_0_d_out_dcbz, loadstore1_0_d_out_load, loadstore1_0_d_out_hold, loadstore1_0_d_out_valid};
  assign n1288_o = dcache_to_loadstore1[0];
  assign n1289_o = dcache_to_loadstore1[64:1];
  assign n1290_o = dcache_to_loadstore1[65];
  assign n1291_o = dcache_to_loadstore1[66];
  assign n1292_o = dcache_to_loadstore1[67];
  assign n1293_o = {loadstore1_0_m_out_rs, loadstore1_0_m_out_addr, loadstore1_0_m_out_sprn, loadstore1_0_m_out_priv, loadstore1_0_m_out_load, loadstore1_0_m_out_iside, loadstore1_0_m_out_mtspr, loadstore1_0_m_out_slbia, loadstore1_0_m_out_tlbie, loadstore1_0_m_out_valid};
  assign n1295_o = mmu_to_loadstore1[0];
  assign n1296_o = mmu_to_loadstore1[1];
  assign n1297_o = mmu_to_loadstore1[2];
  assign n1298_o = mmu_to_loadstore1[3];
  assign n1299_o = mmu_to_loadstore1[4];
  assign n1300_o = mmu_to_loadstore1[5];
  assign n1301_o = mmu_to_loadstore1[6];
  assign n1302_o = mmu_to_loadstore1[70:7];
  assign n1303_o = {loadstore1_0_events_itlb_miss, loadstore1_0_events_store_complete, loadstore1_0_events_load_complete};
  /* core.vhdl:413:5  */
  mmu mmu_0 (
    .clk(clk),
    .rst(core_rst),
    .l_in_valid(n1306_o),
    .l_in_tlbie(n1307_o),
    .l_in_slbia(n1308_o),
    .l_in_mtspr(n1309_o),
    .l_in_iside(n1310_o),
    .l_in_load(n1311_o),
    .l_in_priv(n1312_o),
    .l_in_sprn(n1313_o),
    .l_in_addr(n1314_o),
    .l_in_rs(n1315_o),
    .d_in_stall(n1320_o),
    .d_in_done(n1321_o),
    .d_in_err(n1322_o),
    .d_in_data(n1323_o),
    .l_out_done(mmu_0_l_out_done),
    .l_out_err(mmu_0_l_out_err),
    .l_out_invalid(mmu_0_l_out_invalid),
    .l_out_badtree(mmu_0_l_out_badtree),
    .l_out_segerr(mmu_0_l_out_segerr),
    .l_out_perm_error(mmu_0_l_out_perm_error),
    .l_out_rc_error(mmu_0_l_out_rc_error),
    .l_out_sprval(mmu_0_l_out_sprval),
    .d_out_valid(mmu_0_d_out_valid),
    .d_out_tlbie(mmu_0_d_out_tlbie),
    .d_out_doall(mmu_0_d_out_doall),
    .d_out_tlbld(mmu_0_d_out_tlbld),
    .d_out_addr(mmu_0_d_out_addr),
    .d_out_pte(mmu_0_d_out_pte),
    .i_out_tlbld(mmu_0_i_out_tlbld),
    .i_out_tlbie(mmu_0_i_out_tlbie),
    .i_out_doall(mmu_0_i_out_doall),
    .i_out_addr(mmu_0_i_out_addr),
    .i_out_pte(mmu_0_i_out_pte));
  assign n1306_o = loadstore1_to_mmu[0];
  assign n1307_o = loadstore1_to_mmu[1];
  assign n1308_o = loadstore1_to_mmu[2];
  assign n1309_o = loadstore1_to_mmu[3];
  assign n1310_o = loadstore1_to_mmu[4];
  assign n1311_o = loadstore1_to_mmu[5];
  assign n1312_o = loadstore1_to_mmu[6];
  assign n1313_o = loadstore1_to_mmu[16:7];
  assign n1314_o = loadstore1_to_mmu[80:17];
  assign n1315_o = loadstore1_to_mmu[144:81];
  assign n1316_o = {mmu_0_l_out_sprval, mmu_0_l_out_rc_error, mmu_0_l_out_perm_error, mmu_0_l_out_segerr, mmu_0_l_out_badtree, mmu_0_l_out_invalid, mmu_0_l_out_err, mmu_0_l_out_done};
  assign n1318_o = {mmu_0_d_out_pte, mmu_0_d_out_addr, mmu_0_d_out_tlbld, mmu_0_d_out_doall, mmu_0_d_out_tlbie, mmu_0_d_out_valid};
  assign n1320_o = dcache_to_mmu[0];
  assign n1321_o = dcache_to_mmu[1];
  assign n1322_o = dcache_to_mmu[2];
  assign n1323_o = dcache_to_mmu[66:3];
  assign n1324_o = {mmu_0_i_out_pte, mmu_0_i_out_addr, mmu_0_i_out_doall, mmu_0_i_out_tlbie, mmu_0_i_out_tlbld};
  /* core.vhdl:424:5  */
  dcache_64_4_1_2_2_12_0 dcache_0 (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(clk),
    .rst(rst_dcache),
    .d_in_valid(n1326_o),
    .d_in_hold(n1327_o),
    .d_in_load(n1328_o),
    .d_in_dcbz(n1329_o),
    .d_in_nc(n1330_o),
    .d_in_reserve(n1331_o),
    .d_in_atomic(n1332_o),
    .d_in_atomic_last(n1333_o),
    .d_in_virt_mode(n1334_o),
    .d_in_priv_mode(n1335_o),
    .d_in_addr(n1336_o),
    .d_in_data(n1337_o),
    .d_in_byte_sel(n1338_o),
    .m_in_valid(n1341_o),
    .m_in_tlbie(n1342_o),
    .m_in_doall(n1343_o),
    .m_in_tlbld(n1344_o),
    .m_in_addr(n1345_o),
    .m_in_pte(n1346_o),
    .snoop_in_adr(n1349_o),
    .snoop_in_dat(n1350_o),
    .snoop_in_sel(n1351_o),
    .snoop_in_cyc(n1352_o),
    .snoop_in_stb(n1353_o),
    .snoop_in_we(n1354_o),
    .wishbone_in_dat(n1358_o),
    .wishbone_in_ack(n1359_o),
    .wishbone_in_stall(n1360_o),
    .d_out_valid(dcache_0_d_out_valid),
    .d_out_data(dcache_0_d_out_data),
    .d_out_store_done(dcache_0_d_out_store_done),
    .d_out_error(dcache_0_d_out_error),
    .d_out_cache_paradox(dcache_0_d_out_cache_paradox),
    .m_out_stall(dcache_0_m_out_stall),
    .m_out_done(dcache_0_m_out_done),
    .m_out_err(dcache_0_m_out_err),
    .m_out_data(dcache_0_m_out_data),
    .stall_out(dcache_0_stall_out),
    .wishbone_out_adr(dcache_0_wishbone_out_adr),
    .wishbone_out_dat(dcache_0_wishbone_out_dat),
    .wishbone_out_sel(dcache_0_wishbone_out_sel),
    .wishbone_out_cyc(dcache_0_wishbone_out_cyc),
    .wishbone_out_stb(dcache_0_wishbone_out_stb),
    .wishbone_out_we(dcache_0_wishbone_out_we),
    .events_load_miss(dcache_0_events_load_miss),
    .events_store_miss(dcache_0_events_store_miss),
    .events_dcache_refill(dcache_0_events_dcache_refill),
    .events_dtlb_miss(dcache_0_events_dtlb_miss),
    .events_dtlb_miss_resolved(dcache_0_events_dtlb_miss_resolved),
    .log_out(dcache_0_log_out));
  assign n1326_o = loadstore1_to_dcache[0];
  assign n1327_o = loadstore1_to_dcache[1];
  assign n1328_o = loadstore1_to_dcache[2];
  assign n1329_o = loadstore1_to_dcache[3];
  assign n1330_o = loadstore1_to_dcache[4];
  assign n1331_o = loadstore1_to_dcache[5];
  assign n1332_o = loadstore1_to_dcache[6];
  assign n1333_o = loadstore1_to_dcache[7];
  assign n1334_o = loadstore1_to_dcache[8];
  assign n1335_o = loadstore1_to_dcache[9];
  assign n1336_o = loadstore1_to_dcache[73:10];
  assign n1337_o = loadstore1_to_dcache[137:74];
  assign n1338_o = loadstore1_to_dcache[145:138];
  assign n1339_o = {dcache_0_d_out_cache_paradox, dcache_0_d_out_error, dcache_0_d_out_store_done, dcache_0_d_out_data, dcache_0_d_out_valid};
  assign n1341_o = mmu_to_dcache[0];
  assign n1342_o = mmu_to_dcache[1];
  assign n1343_o = mmu_to_dcache[2];
  assign n1344_o = mmu_to_dcache[3];
  assign n1345_o = mmu_to_dcache[67:4];
  assign n1346_o = mmu_to_dcache[131:68];
  assign n1347_o = {dcache_0_m_out_data, dcache_0_m_out_err, dcache_0_m_out_done, dcache_0_m_out_stall};
  assign n1349_o = n1020_o[28:0];
  assign n1350_o = n1020_o[92:29];
  assign n1351_o = n1020_o[100:93];
  assign n1352_o = n1020_o[101];
  assign n1353_o = n1020_o[102];
  assign n1354_o = n1020_o[103];
  assign n1356_o = {dcache_0_wishbone_out_we, dcache_0_wishbone_out_stb, dcache_0_wishbone_out_cyc, dcache_0_wishbone_out_sel, dcache_0_wishbone_out_dat, dcache_0_wishbone_out_adr};
  assign n1358_o = n1012_o[63:0];
  assign n1359_o = n1012_o[64];
  assign n1360_o = n1012_o[65];
  assign n1361_o = {dcache_0_events_dtlb_miss_resolved, dcache_0_events_dtlb_miss, dcache_0_events_dcache_refill, dcache_0_events_store_miss, dcache_0_events_load_miss};
  /* core.vhdl:448:5  */
  writeback writeback_0 (
    .clk(clk),
    .rst(rst_wback),
    .e_in_valid(n1364_o),
    .e_in_instr_tag(n1365_o),
    .e_in_rc(n1366_o),
    .e_in_mode_32bit(n1367_o),
    .e_in_write_enable(n1368_o),
    .e_in_write_reg(n1369_o),
    .e_in_write_data(n1370_o),
    .e_in_write_cr_enable(n1371_o),
    .e_in_write_cr_mask(n1372_o),
    .e_in_write_cr_data(n1373_o),
    .e_in_write_xerc_enable(n1374_o),
    .e_in_xerc(n1375_o),
    .e_in_interrupt(n1376_o),
    .e_in_intr_vec(n1377_o),
    .e_in_redirect(n1378_o),
    .e_in_redir_mode(n1379_o),
    .e_in_last_nia(n1380_o),
    .e_in_br_offset(n1381_o),
    .e_in_br_last(n1382_o),
    .e_in_br_taken(n1383_o),
    .e_in_abs_br(n1384_o),
    .e_in_srr1(n1385_o),
    .e_in_msr(n1386_o),
    .l_in_valid(n1387_o),
    .l_in_instr_tag(n1388_o),
    .l_in_write_enable(n1389_o),
    .l_in_write_reg(n1390_o),
    .l_in_write_data(n1391_o),
    .l_in_xerc(n1392_o),
    .l_in_rc(n1393_o),
    .l_in_store_done(n1394_o),
    .l_in_interrupt(n1395_o),
    .l_in_intr_vec(n1396_o),
    .l_in_srr0(n1397_o),
    .l_in_srr1(n1398_o),
    .fp_in_valid(n1399_o),
    .fp_in_interrupt(n1400_o),
    .fp_in_instr_tag(n1401_o),
    .fp_in_write_enable(n1402_o),
    .fp_in_write_reg(n1403_o),
    .fp_in_write_data(n1404_o),
    .fp_in_write_cr_enable(n1405_o),
    .fp_in_write_cr_mask(n1406_o),
    .fp_in_write_cr_data(n1407_o),
    .fp_in_intr_vec(n1408_o),
    .fp_in_srr0(n1409_o),
    .fp_in_srr1(n1410_o),
    .w_out_write_reg(writeback_0_w_out_write_reg),
    .w_out_write_data(writeback_0_w_out_write_data),
    .w_out_write_enable(writeback_0_w_out_write_enable),
    .c_out_write_cr_enable(writeback_0_c_out_write_cr_enable),
    .c_out_write_cr_mask(writeback_0_c_out_write_cr_mask),
    .c_out_write_cr_data(writeback_0_c_out_write_cr_data),
    .c_out_write_xerc_enable(writeback_0_c_out_write_xerc_enable),
    .c_out_write_xerc_data(writeback_0_c_out_write_xerc_data),
    .f_out_redirect(writeback_0_f_out_redirect),
    .f_out_virt_mode(writeback_0_f_out_virt_mode),
    .f_out_priv_mode(writeback_0_f_out_priv_mode),
    .f_out_big_endian(writeback_0_f_out_big_endian),
    .f_out_mode_32bit(writeback_0_f_out_mode_32bit),
    .f_out_redirect_nia(writeback_0_f_out_redirect_nia),
    .f_out_br_nia(writeback_0_f_out_br_nia),
    .f_out_br_last(writeback_0_f_out_br_last),
    .f_out_br_taken(writeback_0_f_out_br_taken),
    .events_instr_complete(writeback_0_events_instr_complete),
    .events_fp_complete(writeback_0_events_fp_complete),
    .flush_out(writeback_0_flush_out),
    .interrupt_out(writeback_0_interrupt_out),
    .complete_out_tag(writeback_0_complete_out_tag),
    .complete_out_valid(writeback_0_complete_out_valid));
  assign n1364_o = execute1_to_writeback[0];
  assign n1365_o = execute1_to_writeback[3:1];
  assign n1366_o = execute1_to_writeback[4];
  assign n1367_o = execute1_to_writeback[5];
  assign n1368_o = execute1_to_writeback[6];
  assign n1369_o = execute1_to_writeback[13:7];
  assign n1370_o = execute1_to_writeback[77:14];
  assign n1371_o = execute1_to_writeback[78];
  assign n1372_o = execute1_to_writeback[86:79];
  assign n1373_o = execute1_to_writeback[118:87];
  assign n1374_o = execute1_to_writeback[119];
  assign n1375_o = execute1_to_writeback[124:120];
  assign n1376_o = execute1_to_writeback[125];
  assign n1377_o = execute1_to_writeback[137:126];
  assign n1378_o = execute1_to_writeback[138];
  assign n1379_o = execute1_to_writeback[142:139];
  assign n1380_o = execute1_to_writeback[206:143];
  assign n1381_o = execute1_to_writeback[270:207];
  assign n1382_o = execute1_to_writeback[271];
  assign n1383_o = execute1_to_writeback[272];
  assign n1384_o = execute1_to_writeback[273];
  assign n1385_o = execute1_to_writeback[289:274];
  assign n1386_o = execute1_to_writeback[353:290];
  assign n1387_o = loadstore1_to_writeback[0];
  assign n1388_o = loadstore1_to_writeback[3:1];
  assign n1389_o = loadstore1_to_writeback[4];
  assign n1390_o = loadstore1_to_writeback[11:5];
  assign n1391_o = loadstore1_to_writeback[75:12];
  assign n1392_o = loadstore1_to_writeback[80:76];
  assign n1393_o = loadstore1_to_writeback[81];
  assign n1394_o = loadstore1_to_writeback[82];
  assign n1395_o = loadstore1_to_writeback[83];
  assign n1396_o = loadstore1_to_writeback[95:84];
  assign n1397_o = loadstore1_to_writeback[159:96];
  assign n1398_o = loadstore1_to_writeback[175:160];
  assign n1399_o = fpu_to_writeback[0];
  assign n1400_o = fpu_to_writeback[1];
  assign n1401_o = fpu_to_writeback[4:2];
  assign n1402_o = fpu_to_writeback[5];
  assign n1403_o = fpu_to_writeback[12:6];
  assign n1404_o = fpu_to_writeback[76:13];
  assign n1405_o = fpu_to_writeback[77];
  assign n1406_o = fpu_to_writeback[85:78];
  assign n1407_o = fpu_to_writeback[117:86];
  assign n1408_o = fpu_to_writeback[129:118];
  assign n1409_o = fpu_to_writeback[193:130];
  assign n1410_o = fpu_to_writeback[209:194];
  assign n1411_o = {writeback_0_w_out_write_enable, writeback_0_w_out_write_data, writeback_0_w_out_write_reg};
  assign n1413_o = {writeback_0_c_out_write_xerc_data, writeback_0_c_out_write_xerc_enable, writeback_0_c_out_write_cr_data, writeback_0_c_out_write_cr_mask, writeback_0_c_out_write_cr_enable};
  assign n1415_o = {writeback_0_f_out_br_taken, writeback_0_f_out_br_last, writeback_0_f_out_br_nia, writeback_0_f_out_redirect_nia, writeback_0_f_out_mode_32bit, writeback_0_f_out_big_endian, writeback_0_f_out_priv_mode, writeback_0_f_out_virt_mode, writeback_0_f_out_redirect};
  assign n1417_o = {writeback_0_events_fp_complete, writeback_0_events_instr_complete};
  assign n1421_o = {writeback_0_complete_out_valid, writeback_0_complete_out_tag};
  /* core.vhdl:467:5  */
  core_debug_0 debug_0 (
    .clk(clk),
    .rst(rst_dbg),
    .dmi_addr(dmi_addr),
    .dmi_din(dmi_din),
    .dmi_req(dmi_req),
    .dmi_wr(dmi_wr),
    .terminate(terminate),
    .core_stopped(dbg_core_is_stopped),
    .nia(n1430_o),
    .msr(msr),
    .dbg_gpr_ack(dbg_gpr_ack),
    .dbg_gpr_data(dbg_gpr_data),
    .log_data(log_data),
    .log_read_addr(log_rd_addr),
    .dmi_dout(debug_0_dmi_dout),
    .dmi_ack(debug_0_dmi_ack),
    .core_stop(debug_0_core_stop),
    .core_rst(debug_0_core_rst),
    .icache_rst(debug_0_icache_rst),
    .dbg_gpr_req(debug_0_dbg_gpr_req),
    .dbg_gpr_addr(debug_0_dbg_gpr_addr),
    .log_read_data(debug_0_log_read_data),
    .log_write_addr(debug_0_log_write_addr),
    .terminated_out(debug_0_terminated_out));
  /* core.vhdl:485:37  */
  assign n1430_o = fetch1_to_icache[70:7];
  /* core.vhdl:193:9  */
  always @(posedge clk)
    n1437_q <= core_rst;
  initial
    n1437_q = 1'b1;
  /* core.vhdl:193:9  */
  always @(posedge clk)
    n1439_q <= core_rst;
  initial
    n1439_q = 1'b1;
  /* core.vhdl:193:9  */
  always @(posedge clk)
    n1440_q <= core_rst;
  initial
    n1440_q = 1'b1;
  /* core.vhdl:193:9  */
  always @(posedge clk)
    n1441_q <= core_rst;
  initial
    n1441_q = 1'b1;
  /* core.vhdl:193:9  */
  always @(posedge clk)
    n1442_q <= core_rst;
  initial
    n1442_q = 1'b1;
  /* core.vhdl:193:9  */
  always @(posedge clk)
    n1443_q <= core_rst;
  initial
    n1443_q = 1'b1;
  /* core.vhdl:193:9  */
  always @(posedge clk)
    n1444_q <= core_rst;
  initial
    n1444_q = 1'b1;
  /* core.vhdl:193:9  */
  always @(posedge clk)
    n1445_q <= core_rst;
  initial
    n1445_q = 1'b1;
  /* core.vhdl:193:9  */
  always @(posedge clk)
    n1446_q <= core_rst;
  initial
    n1446_q = 1'b1;
  /* core.vhdl:193:9  */
  always @(posedge clk)
    n1447_q <= rst;
  initial
    n1447_q = 1'b1;
  /* core.vhdl:193:9  */
  always @(posedge clk)
    n1448_q <= alt_reset;
  /* core.vhdl:193:9  */
  assign n1449_o = {register_file_0_log_out, cr_file_0_log_out, dcache_0_log_out, 1'b0, loadstore1_0_log_out, 5'b00000, execute1_0_log_out, decode2_0_log_out, decode1_0_log_out, icache_0_log_out, fetch1_0_log_out};
endmodule

module soc_4096_100000000_0_0_4_0_4_0_4_1_4_4_1_2_2_32_529beb193518cdd5546a21170d32ebafc9f9cb89
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  rst,
   input  system_clk,
   input  [63:0] wb_dram_out_dat,
   input  wb_dram_out_ack,
   input  wb_dram_out_stall,
   input  [31:0] wb_ext_io_out_dat,
   input  wb_ext_io_out_ack,
   input  wb_ext_io_out_stall,
   input  [29:0] wishbone_dma_out_adr,
   input  [31:0] wishbone_dma_out_dat,
   input  [3:0] wishbone_dma_out_sel,
   input  wishbone_dma_out_cyc,
   input  wishbone_dma_out_stb,
   input  wishbone_dma_out_we,
   input  ext_irq_eth,
   input  ext_irq_sdcard,
   input  uart0_rxd,
   input  uart1_rxd,
   input  [3:0] spi_flash_sdat_i,
   input  [31:0] gpio_in,
   input  jtag_tck,
   input  jtag_tdi,
   input  jtag_tms,
   input  jtag_trst,
   input  alt_reset,
   output [28:0] wb_dram_in_adr,
   output [63:0] wb_dram_in_dat,
   output [7:0] wb_dram_in_sel,
   output wb_dram_in_cyc,
   output wb_dram_in_stb,
   output wb_dram_in_we,
   output [29:0] wb_ext_io_in_adr,
   output [31:0] wb_ext_io_in_dat,
   output [3:0] wb_ext_io_in_sel,
   output wb_ext_io_in_cyc,
   output wb_ext_io_in_stb,
   output wb_ext_io_in_we,
   output wb_ext_is_dram_csr,
   output wb_ext_is_dram_init,
   output wb_ext_is_eth,
   output wb_ext_is_sdcard,
   output [31:0] wishbone_dma_in_dat,
   output wishbone_dma_in_ack,
   output wishbone_dma_in_stall,
   output uart0_txd,
   output uart1_txd,
   output spi_flash_sck,
   output spi_flash_cs_n,
   output [3:0] spi_flash_sdat_o,
   output [3:0] spi_flash_sdat_oe,
   output [31:0] gpio_out,
   output [31:0] gpio_dir,
   output jtag_tdo);
  wire [28:0] n71_o;
  wire [63:0] n72_o;
  wire [7:0] n73_o;
  wire n74_o;
  wire n75_o;
  wire n76_o;
  wire [65:0] n77_o;
  wire [29:0] n79_o;
  wire [31:0] n80_o;
  wire [3:0] n81_o;
  wire n82_o;
  wire n83_o;
  wire n84_o;
  wire [33:0] n85_o;
  wire [31:0] n92_o;
  wire n93_o;
  wire n94_o;
  wire [68:0] n95_o;
  wire [65:0] wishbone_dcore_in;
  wire [103:0] wishbone_dcore_out;
  wire [65:0] wishbone_icore_in;
  wire [103:0] wishbone_icore_out;
  wire [65:0] wishbone_debug_in;
  wire [103:0] wishbone_debug_out;
  wire [415:0] wb_masters_out;
  wire [263:0] wb_masters_in;
  wire [65:0] wb_master_in;
  wire [103:0] wb_master_out;
  wire [103:0] wb_snoop;
  wire [103:0] wb_io_in;
  wire [65:0] wb_io_out;
  wire [68:0] wb_sio_out;
  wire [33:0] wb_sio_in;
  wire dram_at_0;
  wire do_core_reset;
  wire [68:0] wb_syscon_in;
  wire [33:0] wb_syscon_out;
  wire [68:0] wb_uart0_in;
  wire [33:0] wb_uart0_out;
  wire [7:0] uart0_dat8;
  wire uart0_irq;
  wire [68:0] wb_uart1_in;
  wire [33:0] wb_uart1_out;
  wire uart1_irq;
  wire [68:0] wb_spiflash_in;
  wire [33:0] wb_spiflash_out;
  wire wb_spiflash_is_reg;
  wire wb_spiflash_is_map;
  wire [68:0] wb_xics_icp_in;
  wire [33:0] wb_xics_icp_out;
  wire [68:0] wb_xics_ics_in;
  wire [33:0] wb_xics_ics_out;
  wire [15:0] int_level_in;
  wire [11:0] ics_to_icp;
  wire core_ext_irq;
  wire [68:0] wb_gpio_in;
  wire [33:0] wb_gpio_out;
  reg gpio_intr;
  wire [103:0] wb_bram_in;
  wire [65:0] wb_bram_out;
  wire [7:0] dmi_addr;
  wire [63:0] dmi_din;
  wire [63:0] dmi_dout;
  wire dmi_req;
  wire dmi_wr;
  wire dmi_ack;
  wire [63:0] dmi_wb_dout;
  wire dmi_wb_req;
  wire dmi_wb_ack;
  wire [63:0] dmi_core_dout;
  wire dmi_core_req;
  wire dmi_core_ack;
  reg rst_core;
  reg rst_uart;
  reg rst_xics;
  reg rst_spi;
  reg rst_gpio;
  reg rst_bram;
  reg rst_dtm;
  reg rst_wbar;
  reg rst_wbdb;
  wire alt_reset_d;
  wire [2:0] current_io_decode;
  wire io_cycle_none;
  wire io_cycle_syscon;
  wire io_cycle_uart;
  wire io_cycle_uart1;
  wire io_cycle_icp;
  wire io_cycle_ics;
  wire io_cycle_spi_flash;
  wire io_cycle_gpio;
  wire io_cycle_external;
  wire n117_o;
  wire [28:0] processor_wishbone_insn_out_adr;
  wire [63:0] processor_wishbone_insn_out_dat;
  wire [7:0] processor_wishbone_insn_out_sel;
  wire processor_wishbone_insn_out_cyc;
  wire processor_wishbone_insn_out_stb;
  wire processor_wishbone_insn_out_we;
  wire [28:0] processor_wishbone_data_out_adr;
  wire [63:0] processor_wishbone_data_out_dat;
  wire [7:0] processor_wishbone_data_out_sel;
  wire processor_wishbone_data_out_cyc;
  wire processor_wishbone_data_out_stb;
  wire processor_wishbone_data_out_we;
  wire [63:0] processor_dmi_dout;
  wire processor_dmi_ack;
  wire processor_terminated_out;
  wire [63:0] n129_o;
  wire n130_o;
  wire n131_o;
  wire [103:0] n132_o;
  wire [63:0] n134_o;
  wire n135_o;
  wire n136_o;
  wire [103:0] n137_o;
  wire [28:0] n139_o;
  wire [63:0] n140_o;
  wire [7:0] n141_o;
  wire n142_o;
  wire n143_o;
  wire n144_o;
  wire [3:0] n145_o;
  wire [28:0] n154_o;
  wire [31:0] n157_o;
  wire [31:0] n158_o;
  wire [63:0] n159_o;
  localparam [7:0] n161_o = 8'b00000000;
  wire n163_o;
  wire n164_o;
  wire [3:0] n165_o;
  wire [3:0] n166_o;
  wire [3:0] n167_o;
  wire [3:0] n168_o;
  wire [3:0] n169_o;
  wire [3:0] n170_o;
  wire n172_o;
  wire n174_o;
  wire n176_o;
  wire [103:0] n177_o;
  wire [415:0] n178_o;
  wire [65:0] n179_o;
  wire [65:0] n180_o;
  wire [65:0] n182_o;
  wire [29:0] n183_o;
  wire n189_o;
  wire n193_o;
  wire n194_o;
  wire n195_o;
  wire [31:0] n196_o;
  wire [31:0] n197_o;
  wire [31:0] n198_o;
  wire [33:0] n199_o;
  wire [65:0] n200_o;
  wire [263:0] wishbone_arbiter_0_wb_masters_out;
  wire [28:0] wishbone_arbiter_0_wb_slave_out_adr;
  wire [63:0] wishbone_arbiter_0_wb_slave_out_dat;
  wire [7:0] wishbone_arbiter_0_wb_slave_out_sel;
  wire wishbone_arbiter_0_wb_slave_out_cyc;
  wire wishbone_arbiter_0_wb_slave_out_stb;
  wire wishbone_arbiter_0_wb_slave_out_we;
  wire [103:0] n202_o;
  wire [63:0] n204_o;
  wire n205_o;
  wire n206_o;
  wire n209_o;
  wire n211_o;
  wire n212_o;
  wire n213_o;
  wire [101:0] n214_o;
  wire [2:0] n219_o;
  wire [3:0] n220_o;
  wire [3:0] n223_o;
  wire n224_o;
  wire [3:0] n227_o;
  wire n228_o;
  wire [3:0] n231_o;
  wire n232_o;
  wire [3:0] n235_o;
  wire n236_o;
  wire [3:0] n239_o;
  wire n240_o;
  wire [1:0] n243_o;
  wire [1:0] n245_o;
  wire [1:0] n247_o;
  wire [1:0] n249_o;
  wire [1:0] n251_o;
  wire [1:0] n254_o;
  wire [100:0] n255_o;
  wire [1:0] n257_o;
  wire [100:0] n258_o;
  wire [1:0] n260_o;
  wire [100:0] n261_o;
  wire n262_o;
  wire n264_o;
  wire n265_o;
  wire n267_o;
  wire n268_o;
  wire n270_o;
  wire [2:0] n271_o;
  reg n273_o;
  reg [65:0] n275_o;
  reg n277_o;
  reg n279_o;
  reg [1:0] slave_io_latch_state;
  reg slave_io_latch_has_top;
  wire n294_o;
  wire n295_o;
  wire n296_o;
  wire n299_o;
  wire [28:0] n300_o;
  wire [29:0] n302_o;
  wire [3:0] n303_o;
  wire n305_o;
  wire [3:0] n306_o;
  wire n308_o;
  wire n309_o;
  wire [31:0] n310_o;
  wire [31:0] n311_o;
  wire [31:0] n312_o;
  wire [3:0] n313_o;
  wire n314_o;
  wire [31:0] n315_o;
  wire [31:0] n316_o;
  wire [31:0] n317_o;
  wire [3:0] n318_o;
  wire [35:0] n320_o;
  wire [35:0] n321_o;
  wire n322_o;
  wire n323_o;
  wire [35:0] n324_o;
  wire [28:0] n325_o;
  wire [1:0] n328_o;
  wire n329_o;
  wire n330_o;
  wire [65:0] n331_o;
  wire [1:0] n332_o;
  wire [65:0] n333_o;
  wire [65:0] n334_o;
  wire [1:0] n335_o;
  wire [1:0] n336_o;
  wire [1:0] n337_o;
  wire n338_o;
  wire n342_o;
  wire n344_o;
  wire n345_o;
  wire n346_o;
  wire n348_o;
  wire n349_o;
  wire n350_o;
  wire n351_o;
  wire n352_o;
  wire [31:0] n353_o;
  wire [31:0] n354_o;
  wire [31:0] n355_o;
  wire n356_o;
  wire [31:0] n357_o;
  wire [31:0] n358_o;
  wire [31:0] n359_o;
  wire [3:0] n360_o;
  wire [1:0] n365_o;
  wire [1:0] n366_o;
  wire [1:0] n367_o;
  wire [35:0] n368_o;
  wire n369_o;
  wire n370_o;
  wire [35:0] n371_o;
  wire [35:0] n372_o;
  wire n373_o;
  wire [1:0] n376_o;
  wire n379_o;
  wire n381_o;
  wire [1:0] n382_o;
  wire [1:0] n383_o;
  wire n385_o;
  wire n387_o;
  wire n388_o;
  wire [1:0] n389_o;
  wire n391_o;
  wire n393_o;
  wire n394_o;
  wire n395_o;
  wire n397_o;
  wire n398_o;
  wire n399_o;
  wire n400_o;
  wire n401_o;
  wire [31:0] n402_o;
  wire [31:0] n403_o;
  wire [31:0] n404_o;
  wire [33:0] n407_o;
  wire [33:0] n408_o;
  wire [33:0] n409_o;
  wire [1:0] n411_o;
  wire n414_o;
  wire n416_o;
  wire [2:0] n417_o;
  wire [31:0] n418_o;
  reg [31:0] n420_o;
  wire [31:0] n421_o;
  wire [31:0] n422_o;
  reg [31:0] n424_o;
  wire n425_o;
  wire n426_o;
  reg n428_o;
  wire n429_o;
  wire n430_o;
  reg n432_o;
  wire n433_o;
  wire n434_o;
  reg n436_o;
  wire [28:0] n437_o;
  wire [28:0] n438_o;
  reg [28:0] n440_o;
  wire [35:0] n441_o;
  wire [35:0] n442_o;
  reg [35:0] n444_o;
  wire n445_o;
  reg n447_o;
  wire n448_o;
  wire n449_o;
  reg n451_o;
  reg [1:0] n453_o;
  reg n455_o;
  reg n460_o;
  reg n463_o;
  wire [65:0] n464_o;
  wire [1:0] n465_o;
  wire [63:0] n466_o;
  wire [63:0] n467_o;
  wire [63:0] n468_o;
  wire [1:0] n469_o;
  wire [1:0] n470_o;
  wire [65:0] n471_o;
  wire [1:0] n472_o;
  wire [65:0] n473_o;
  wire [65:0] n474_o;
  wire n475_o;
  wire n476_o;
  wire n477_o;
  wire n478_o;
  wire n479_o;
  wire [1:0] n481_o;
  wire n483_o;
  wire n487_o;
  wire n490_o;
  wire n492_o;
  wire n495_o;
  wire n497_o;
  wire n502_o;
  wire n503_o;
  wire n505_o;
  wire n507_o;
  wire n509_o;
  wire n511_o;
  wire n513_o;
  wire n515_o;
  wire n517_o;
  wire n519_o;
  wire n521_o;
  wire n523_o;
  wire n525_o;
  wire [17:0] n526_o;
  wire [19:0] n528_o;
  wire [19:0] n531_o;
  wire n532_o;
  wire n534_o;
  wire [19:0] n537_o;
  wire n538_o;
  wire [19:0] n541_o;
  wire n542_o;
  wire [19:0] n545_o;
  wire n546_o;
  wire n548_o;
  wire n563_o;
  wire n565_o;
  wire n567_o;
  wire [2:0] n570_o;
  wire [19:0] n573_o;
  wire n574_o;
  wire [19:0] n577_o;
  wire n578_o;
  wire [19:0] n581_o;
  wire n582_o;
  wire [19:0] n585_o;
  wire n586_o;
  wire [19:0] n589_o;
  wire n590_o;
  wire [19:0] n593_o;
  wire n594_o;
  wire [19:0] n597_o;
  wire n598_o;
  wire n600_o;
  wire n602_o;
  wire [2:0] n605_o;
  wire n607_o;
  wire n608_o;
  wire n610_o;
  wire n611_o;
  wire [2:0] n613_o;
  wire n614_o;
  wire n615_o;
  wire n617_o;
  wire n618_o;
  wire n619_o;
  wire [2:0] n621_o;
  wire n622_o;
  wire n623_o;
  wire n625_o;
  wire n626_o;
  wire n627_o;
  wire n628_o;
  wire [2:0] n630_o;
  wire n631_o;
  wire n632_o;
  wire n634_o;
  wire n635_o;
  wire n636_o;
  wire n637_o;
  wire n638_o;
  wire [2:0] n640_o;
  wire n641_o;
  wire n642_o;
  wire n644_o;
  wire n645_o;
  wire n646_o;
  wire n647_o;
  wire n648_o;
  wire n649_o;
  wire [2:0] n651_o;
  wire n652_o;
  wire n653_o;
  wire n655_o;
  wire n656_o;
  wire n657_o;
  wire n658_o;
  wire n659_o;
  wire n660_o;
  wire n661_o;
  wire [2:0] n663_o;
  wire n664_o;
  wire n665_o;
  wire n666_o;
  wire n667_o;
  wire n668_o;
  wire n669_o;
  wire n670_o;
  wire n671_o;
  wire n672_o;
  wire n673_o;
  wire n674_o;
  wire [2:0] n675_o;
  wire n676_o;
  wire n677_o;
  wire n679_o;
  wire n680_o;
  wire n681_o;
  wire n682_o;
  wire n683_o;
  wire n684_o;
  wire n685_o;
  wire n687_o;
  wire n688_o;
  wire n689_o;
  wire [2:0] n691_o;
  wire n692_o;
  wire n694_o;
  wire n695_o;
  wire n696_o;
  wire n697_o;
  wire n698_o;
  wire n699_o;
  wire n700_o;
  wire n701_o;
  wire n702_o;
  wire n703_o;
  wire n704_o;
  wire n706_o;
  wire [2:0] n708_o;
  wire n711_o;
  wire n712_o;
  wire n713_o;
  wire n714_o;
  wire n715_o;
  wire n717_o;
  wire n718_o;
  wire n719_o;
  wire n720_o;
  wire n721_o;
  wire n722_o;
  wire n723_o;
  wire n724_o;
  wire n725_o;
  wire [65:0] n732_o;
  wire [68:0] n734_o;
  reg [1:0] n756_q;
  reg n757_q;
  wire [1:0] n760_o;
  wire [65:0] n761_o;
  wire [1:0] n762_o;
  wire [65:0] n763_o;
  wire [1:0] n764_o;
  wire [37:0] n767_o;
  wire [25:0] n768_o;
  wire [1:0] n769_o;
  wire [65:0] n770_o;
  localparam [29:0] n771_o = 30'b000000000000000000000000000000;
  wire [5:0] n773_o;
  wire [23:0] n774_o;
  wire [1:0] n775_o;
  wire [35:0] n776_o;
  localparam [29:0] n777_o = 30'b000000000000000000000000000000;
  wire [9:0] n779_o;
  wire [19:0] n780_o;
  wire [1:0] n781_o;
  wire [35:0] n782_o;
  wire [1:0] n783_o;
  wire [65:0] n784_o;
  wire [1:0] n785_o;
  wire [65:0] n786_o;
  wire n788_o;
  wire n790_o;
  wire n792_o;
  wire n794_o;
  wire n796_o;
  wire n798_o;
  wire n800_o;
  wire n802_o;
  wire [7:0] n803_o;
  reg [33:0] n805_o;
  wire n807_o;
  wire n808_o;
  wire n809_o;
  wire [33:0] n811_o;
  wire [33:0] n812_o;
  wire [31:0] syscon0_wishbone_out_dat;
  wire syscon0_wishbone_out_ack;
  wire syscon0_wishbone_out_stall;
  wire syscon0_dram_at_0;
  wire syscon0_core_reset;
  wire syscon0_soc_reset;
  wire [29:0] n814_o;
  wire [31:0] n815_o;
  wire [3:0] n816_o;
  wire n817_o;
  wire n818_o;
  wire n819_o;
  wire [33:0] n820_o;
  wire uart0_16550_irq_l;
  wire [7:0] uart0_16550_uart0_wb_dat_o;
  wire uart0_16550_uart0_wb_ack_o;
  wire uart0_16550_uart0_int_o;
  wire uart0_16550_uart0_stx_pad_o;
  wire uart0_16550_uart0_rts_pad_o;
  wire uart0_16550_uart0_dtr_pad_o;
  wire [2:0] n824_o;
  wire [7:0] n825_o;
  wire n827_o;
  wire n828_o;
  wire n829_o;
  localparam n833_o = 1'b1;
  localparam n834_o = 1'b1;
  localparam n835_o = 1'b0;
  localparam n836_o = 1'b1;
  wire [31:0] n842_o;
  wire n843_o;
  wire n844_o;
  wire n846_o;
  wire n847_o;
  wire n848_o;
  wire [31:0] spiflash_gen_spiflash_wb_out_dat;
  wire spiflash_gen_spiflash_wb_out_ack;
  wire spiflash_gen_spiflash_wb_out_stall;
  wire spiflash_gen_spiflash_sck;
  wire spiflash_gen_spiflash_cs_n;
  wire [3:0] spiflash_gen_spiflash_sdat_o;
  wire [3:0] spiflash_gen_spiflash_sdat_oe;
  wire [29:0] n851_o;
  wire [31:0] n852_o;
  wire [3:0] n853_o;
  wire n854_o;
  wire n855_o;
  wire n856_o;
  wire [33:0] n857_o;
  wire [31:0] xics_icp_wb_out_dat;
  wire xics_icp_wb_out_ack;
  wire xics_icp_wb_out_stall;
  wire xics_icp_core_irq_out;
  wire [29:0] n863_o;
  wire [31:0] n864_o;
  wire [3:0] n865_o;
  wire n866_o;
  wire n867_o;
  wire n868_o;
  wire [33:0] n869_o;
  wire [3:0] n871_o;
  wire [7:0] n872_o;
  wire [31:0] xics_ics_wb_out_dat;
  wire xics_ics_wb_out_ack;
  wire xics_ics_wb_out_stall;
  wire [3:0] xics_ics_icp_out_src;
  wire [7:0] xics_ics_icp_out_pri;
  wire [29:0] n874_o;
  wire [31:0] n875_o;
  wire [3:0] n876_o;
  wire n877_o;
  wire n878_o;
  wire n879_o;
  wire [33:0] n880_o;
  wire [11:0] n882_o;
  wire [31:0] gpio0_gen_gpio_wb_out_dat;
  wire gpio0_gen_gpio_wb_out_ack;
  wire gpio0_gen_gpio_wb_out_stall;
  wire [31:0] gpio0_gen_gpio_gpio_out;
  wire [31:0] gpio0_gen_gpio_gpio_dir;
  wire gpio0_gen_gpio_intr;
  wire [29:0] n884_o;
  wire [31:0] n885_o;
  wire [3:0] n886_o;
  wire n887_o;
  wire n888_o;
  wire n889_o;
  wire [33:0] n890_o;
  localparam [15:0] n896_o = 16'b0000000000000000;
  wire [10:0] n901_o;
  wire [63:0] bram_bram0_wishbone_out_dat;
  wire bram_bram0_wishbone_out_ack;
  wire bram_bram0_wishbone_out_stall;
  wire [28:0] n903_o;
  wire [63:0] n904_o;
  wire [7:0] n905_o;
  wire n906_o;
  wire n907_o;
  wire n908_o;
  wire [65:0] n909_o;
  wire [7:0] dmi_jtag_dtm_dmi_addr;
  wire [63:0] dmi_jtag_dtm_dmi_dout;
  wire dmi_jtag_dtm_dmi_req;
  wire dmi_jtag_dtm_dmi_wr;
  wire dmi_jtag_dtm_jtag_tdo;
  wire [7:0] n920_o;
  wire n921_o;
  wire [7:0] n924_o;
  wire n925_o;
  wire [1:0] n928_o;
  wire [1:0] n930_o;
  wire n933_o;
  wire n935_o;
  wire [1:0] n936_o;
  reg [63:0] n938_o;
  reg n939_o;
  reg n941_o;
  reg n944_o;
  wire [63:0] wishbone_debug_dmi_dout;
  wire wishbone_debug_dmi_ack;
  wire [28:0] wishbone_debug_wb_out_adr;
  wire [63:0] wishbone_debug_wb_out_dat;
  wire [7:0] wishbone_debug_wb_out_sel;
  wire wishbone_debug_wb_out_cyc;
  wire wishbone_debug_wb_out_stb;
  wire wishbone_debug_wb_out_we;
  wire [1:0] n947_o;
  wire [103:0] n950_o;
  wire [63:0] n952_o;
  wire n953_o;
  wire n954_o;
  wire [103:0] n955_o;
  wire [103:0] n956_o;
  reg [65:0] n957_q;
  reg [68:0] n958_q;
  wire [68:0] n959_o;
  wire [68:0] n960_o;
  wire [33:0] n961_o;
  reg n962_q;
  wire [68:0] n963_o;
  wire [33:0] n964_o;
  wire [68:0] n966_o;
  reg n967_q;
  reg n968_q;
  wire [68:0] n969_o;
  wire [68:0] n970_o;
  wire [15:0] n971_o;
  wire [68:0] n972_o;
  wire [103:0] n973_o;
  reg n974_q;
  reg n975_q;
  reg n976_q;
  reg n977_q;
  reg n978_q;
  reg n979_q;
  reg n980_q;
  reg n981_q;
  reg n982_q;
  reg n983_q;
  wire [2:0] n984_o;
  reg [2:0] n985_q;
  reg n986_q;
  reg n987_q;
  reg n988_q;
  reg n989_q;
  reg n990_q;
  reg n991_q;
  reg n992_q;
  reg n993_q;
  reg n994_q;
  wire [103:0] n995_o;
  wire [68:0] n996_o;
  reg n997_q;
  reg n998_q;
  wire n999_o;
  reg n1000_q;
  wire n1001_o;
  reg n1002_q;
  localparam n1003_o = 1'bZ;
  assign wb_dram_in_adr = n71_o;
  assign wb_dram_in_dat = n72_o;
  assign wb_dram_in_sel = n73_o;
  assign wb_dram_in_cyc = n74_o;
  assign wb_dram_in_stb = n75_o;
  assign wb_dram_in_we = n76_o;
  assign wb_ext_io_in_adr = n79_o;
  assign wb_ext_io_in_dat = n80_o;
  assign wb_ext_io_in_sel = n81_o;
  assign wb_ext_io_in_cyc = n82_o;
  assign wb_ext_io_in_stb = n83_o;
  assign wb_ext_io_in_we = n84_o;
  assign wb_ext_is_dram_csr = n997_q;
  assign wb_ext_is_dram_init = n998_q;
  assign wb_ext_is_eth = n1000_q;
  assign wb_ext_is_sdcard = n1002_q;
  assign wishbone_dma_in_dat = n92_o;
  assign wishbone_dma_in_ack = n93_o;
  assign wishbone_dma_in_stall = n94_o;
  assign uart0_txd = uart0_16550_uart0_stx_pad_o;
  assign uart1_txd = n1003_o;
  assign spi_flash_sck = spiflash_gen_spiflash_sck;
  assign spi_flash_cs_n = spiflash_gen_spiflash_cs_n;
  assign spi_flash_sdat_o = spiflash_gen_spiflash_sdat_o;
  assign spi_flash_sdat_oe = spiflash_gen_spiflash_sdat_oe;
  assign gpio_out = gpio0_gen_gpio_gpio_out;
  assign gpio_dir = gpio0_gen_gpio_gpio_dir;
  assign jtag_tdo = dmi_jtag_dtm_jtag_tdo;
  /* asic/top-asic.vhdl:278:34  */
  assign n71_o = n995_o[28:0];
  /* asic/top-asic.vhdl:277:34  */
  assign n72_o = n995_o[92:29];
  /* asic/top-asic.vhdl:275:34  */
  assign n73_o = n995_o[100:93];
  /* asic/top-asic.vhdl:274:34  */
  assign n74_o = n995_o[101];
  /* asic/top-asic.vhdl:273:34  */
  assign n75_o = n995_o[102];
  /* asic/top-asic.vhdl:265:34  */
  assign n76_o = n995_o[103];
  /* asic/top-asic.vhdl:264:34  */
  assign n77_o = {wb_dram_out_stall, wb_dram_out_ack, wb_dram_out_dat};
  /* asic/top-asic.vhdl:211:34  */
  assign n79_o = n996_o[29:0];
  /* asic/top-asic.vhdl:204:34  */
  assign n80_o = n996_o[61:30];
  /* asic/top-asic.vhdl:203:34  */
  assign n81_o = n996_o[65:62];
  /* asic/top-asic.vhdl:198:34  */
  assign n82_o = n996_o[66];
  /* asic/top-asic.vhdl:197:34  */
  assign n83_o = n996_o[67];
  /* asic/top-asic.vhdl:196:34  */
  assign n84_o = n996_o[68];
  /* asic/top-asic.vhdl:195:34  */
  assign n85_o = {wb_ext_io_out_stall, wb_ext_io_out_ack, wb_ext_io_out_dat};
  /* asic/top-asic.vhdl:67:9  */
  assign n92_o = n199_o[31:0];
  /* asic/top-asic.vhdl:66:9  */
  assign n93_o = n199_o[32];
  /* asic/top-asic.vhdl:63:9  */
  assign n94_o = n199_o[33];
  /* asic/top-asic.vhdl:56:9  */
  assign n95_o = {wishbone_dma_out_we, wishbone_dma_out_stb, wishbone_dma_out_cyc, wishbone_dma_out_sel, wishbone_dma_out_dat, wishbone_dma_out_adr};
  /* soc.vhdl:149:12  */
  assign wishbone_dcore_in = n179_o; // (signal)
  /* soc.vhdl:150:12  */
  assign wishbone_dcore_out = n137_o; // (signal)
  /* soc.vhdl:151:12  */
  assign wishbone_icore_in = n180_o; // (signal)
  /* soc.vhdl:152:12  */
  assign wishbone_icore_out = n132_o; // (signal)
  /* soc.vhdl:153:12  */
  assign wishbone_debug_in = n200_o; // (signal)
  /* soc.vhdl:154:12  */
  assign wishbone_debug_out = n950_o; // (signal)
  /* soc.vhdl:159:12  */
  assign wb_masters_out = n178_o; // (signal)
  /* soc.vhdl:160:12  */
  assign wb_masters_in = wishbone_arbiter_0_wb_masters_out; // (signal)
  /* soc.vhdl:163:12  */
  assign wb_master_in = n275_o; // (signal)
  /* soc.vhdl:164:12  */
  assign wb_master_out = n202_o; // (signal)
  /* soc.vhdl:165:12  */
  assign wb_snoop = n955_o; // (signal)
  /* soc.vhdl:168:12  */
  assign wb_io_in = n956_o; // (signal)
  /* soc.vhdl:169:12  */
  assign wb_io_out = n957_q; // (signal)
  /* soc.vhdl:172:12  */
  assign wb_sio_out = n958_q; // (signal)
  /* soc.vhdl:173:12  */
  assign wb_sio_in = n812_o; // (signal)
  /* soc.vhdl:176:12  */
  assign dram_at_0 = syscon0_dram_at_0; // (signal)
  /* soc.vhdl:177:12  */
  assign do_core_reset = syscon0_core_reset; // (signal)
  /* soc.vhdl:178:12  */
  assign wb_syscon_in = n959_o; // (signal)
  /* soc.vhdl:179:12  */
  assign wb_syscon_out = n820_o; // (signal)
  /* soc.vhdl:182:12  */
  assign wb_uart0_in = n960_o; // (signal)
  /* soc.vhdl:183:12  */
  assign wb_uart0_out = n961_o; // (signal)
  /* soc.vhdl:184:12  */
  assign uart0_dat8 = uart0_16550_uart0_wb_dat_o; // (signal)
  /* soc.vhdl:185:12  */
  assign uart0_irq = n962_q; // (signal)
  /* soc.vhdl:188:12  */
  assign wb_uart1_in = n963_o; // (signal)
  /* soc.vhdl:189:12  */
  assign wb_uart1_out = n964_o; // (signal)
  /* soc.vhdl:191:12  */
  assign uart1_irq = 1'b0; // (signal)
  /* soc.vhdl:194:12  */
  assign wb_spiflash_in = n966_o; // (signal)
  /* soc.vhdl:195:12  */
  assign wb_spiflash_out = n857_o; // (signal)
  /* soc.vhdl:196:12  */
  assign wb_spiflash_is_reg = n967_q; // (signal)
  /* soc.vhdl:197:12  */
  assign wb_spiflash_is_map = n968_q; // (signal)
  /* soc.vhdl:200:12  */
  assign wb_xics_icp_in = n969_o; // (signal)
  /* soc.vhdl:201:12  */
  assign wb_xics_icp_out = n869_o; // (signal)
  /* soc.vhdl:202:12  */
  assign wb_xics_ics_in = n970_o; // (signal)
  /* soc.vhdl:203:12  */
  assign wb_xics_ics_out = n880_o; // (signal)
  /* soc.vhdl:204:12  */
  assign int_level_in = n971_o; // (signal)
  /* soc.vhdl:205:12  */
  assign ics_to_icp = n882_o; // (signal)
  /* soc.vhdl:206:12  */
  assign core_ext_irq = xics_icp_core_irq_out; // (signal)
  /* soc.vhdl:209:12  */
  assign wb_gpio_in = n972_o; // (signal)
  /* soc.vhdl:210:12  */
  assign wb_gpio_out = n890_o; // (signal)
  /* soc.vhdl:211:12  */
  always @*
    gpio_intr = gpio0_gen_gpio_intr; // (isignal)
  initial
    gpio_intr = 1'b0;
  /* soc.vhdl:214:12  */
  assign wb_bram_in = n973_o; // (signal)
  /* soc.vhdl:215:12  */
  assign wb_bram_out = n909_o; // (signal)
  /* soc.vhdl:218:12  */
  assign dmi_addr = dmi_jtag_dtm_dmi_addr; // (signal)
  /* soc.vhdl:219:12  */
  assign dmi_din = n938_o; // (signal)
  /* soc.vhdl:220:12  */
  assign dmi_dout = dmi_jtag_dtm_dmi_dout; // (signal)
  /* soc.vhdl:221:12  */
  assign dmi_req = dmi_jtag_dtm_dmi_req; // (signal)
  /* soc.vhdl:222:12  */
  assign dmi_wr = dmi_jtag_dtm_dmi_wr; // (signal)
  /* soc.vhdl:223:12  */
  assign dmi_ack = n939_o; // (signal)
  /* soc.vhdl:226:12  */
  assign dmi_wb_dout = wishbone_debug_dmi_dout; // (signal)
  /* soc.vhdl:227:12  */
  assign dmi_wb_req = n941_o; // (signal)
  /* soc.vhdl:228:12  */
  assign dmi_wb_ack = wishbone_debug_dmi_ack; // (signal)
  /* soc.vhdl:229:12  */
  assign dmi_core_dout = processor_dmi_dout; // (signal)
  /* soc.vhdl:230:12  */
  assign dmi_core_req = n944_o; // (signal)
  /* soc.vhdl:231:12  */
  assign dmi_core_ack = processor_dmi_ack; // (signal)
  /* soc.vhdl:234:12  */
  always @*
    rst_core = n974_q; // (isignal)
  initial
    rst_core = 1'b1;
  /* soc.vhdl:235:12  */
  always @*
    rst_uart = n975_q; // (isignal)
  initial
    rst_uart = 1'b1;
  /* soc.vhdl:236:12  */
  always @*
    rst_xics = n976_q; // (isignal)
  initial
    rst_xics = 1'b1;
  /* soc.vhdl:237:12  */
  always @*
    rst_spi = n977_q; // (isignal)
  initial
    rst_spi = 1'b1;
  /* soc.vhdl:238:12  */
  always @*
    rst_gpio = n978_q; // (isignal)
  initial
    rst_gpio = 1'b1;
  /* soc.vhdl:239:12  */
  always @*
    rst_bram = n979_q; // (isignal)
  initial
    rst_bram = 1'b1;
  /* soc.vhdl:240:12  */
  always @*
    rst_dtm = n980_q; // (isignal)
  initial
    rst_dtm = 1'b1;
  /* soc.vhdl:241:12  */
  always @*
    rst_wbar = n981_q; // (isignal)
  initial
    rst_wbar = 1'b1;
  /* soc.vhdl:242:12  */
  always @*
    rst_wbdb = n982_q; // (isignal)
  initial
    rst_wbdb = 1'b1;
  /* soc.vhdl:243:12  */
  assign alt_reset_d = n983_q; // (signal)
  /* soc.vhdl:254:12  */
  assign current_io_decode = n985_q; // (signal)
  /* soc.vhdl:256:12  */
  assign io_cycle_none = n986_q; // (signal)
  /* soc.vhdl:257:12  */
  assign io_cycle_syscon = n987_q; // (signal)
  /* soc.vhdl:258:12  */
  assign io_cycle_uart = n988_q; // (signal)
  /* soc.vhdl:259:12  */
  assign io_cycle_uart1 = n989_q; // (signal)
  /* soc.vhdl:260:12  */
  assign io_cycle_icp = n990_q; // (signal)
  /* soc.vhdl:261:12  */
  assign io_cycle_ics = n991_q; // (signal)
  /* soc.vhdl:262:12  */
  assign io_cycle_spi_flash = n992_q; // (signal)
  /* soc.vhdl:263:12  */
  assign io_cycle_gpio = n993_q; // (signal)
  /* soc.vhdl:264:12  */
  assign io_cycle_external = n994_q; // (signal)
  /* soc.vhdl:327:32  */
  assign n117_o = rst | do_core_reset;
  /* soc.vhdl:341:5  */
  core_0_4_1_4_4_1_2_2_452bf2882a9b5f1c06340d5059c72dbd8af3bf8b processor (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(system_clk),
    .rst(rst_core),
    .alt_reset(alt_reset_d),
    .wishbone_insn_in_dat(n129_o),
    .wishbone_insn_in_ack(n130_o),
    .wishbone_insn_in_stall(n131_o),
    .wishbone_data_in_dat(n134_o),
    .wishbone_data_in_ack(n135_o),
    .wishbone_data_in_stall(n136_o),
    .wb_snoop_in_adr(n139_o),
    .wb_snoop_in_dat(n140_o),
    .wb_snoop_in_sel(n141_o),
    .wb_snoop_in_cyc(n142_o),
    .wb_snoop_in_stb(n143_o),
    .wb_snoop_in_we(n144_o),
    .dmi_addr(n145_o),
    .dmi_din(dmi_dout),
    .dmi_req(dmi_core_req),
    .dmi_wr(dmi_wr),
    .ext_irq(core_ext_irq),
    .wishbone_insn_out_adr(processor_wishbone_insn_out_adr),
    .wishbone_insn_out_dat(processor_wishbone_insn_out_dat),
    .wishbone_insn_out_sel(processor_wishbone_insn_out_sel),
    .wishbone_insn_out_cyc(processor_wishbone_insn_out_cyc),
    .wishbone_insn_out_stb(processor_wishbone_insn_out_stb),
    .wishbone_insn_out_we(processor_wishbone_insn_out_we),
    .wishbone_data_out_adr(processor_wishbone_data_out_adr),
    .wishbone_data_out_dat(processor_wishbone_data_out_dat),
    .wishbone_data_out_sel(processor_wishbone_data_out_sel),
    .wishbone_data_out_cyc(processor_wishbone_data_out_cyc),
    .wishbone_data_out_stb(processor_wishbone_data_out_stb),
    .wishbone_data_out_we(processor_wishbone_data_out_we),
    .dmi_dout(processor_dmi_dout),
    .dmi_ack(processor_dmi_ack),
    .terminated_out());
  assign n129_o = wishbone_icore_in[63:0];
  assign n130_o = wishbone_icore_in[64];
  assign n131_o = wishbone_icore_in[65];
  assign n132_o = {processor_wishbone_insn_out_we, processor_wishbone_insn_out_stb, processor_wishbone_insn_out_cyc, processor_wishbone_insn_out_sel, processor_wishbone_insn_out_dat, processor_wishbone_insn_out_adr};
  assign n134_o = wishbone_dcore_in[63:0];
  assign n135_o = wishbone_dcore_in[64];
  assign n136_o = wishbone_dcore_in[65];
  assign n137_o = {processor_wishbone_data_out_we, processor_wishbone_data_out_stb, processor_wishbone_data_out_cyc, processor_wishbone_data_out_sel, processor_wishbone_data_out_dat, processor_wishbone_data_out_adr};
  assign n139_o = wb_snoop[28:0];
  assign n140_o = wb_snoop[92:29];
  assign n141_o = wb_snoop[100:93];
  assign n142_o = wb_snoop[101];
  assign n143_o = wb_snoop[102];
  assign n144_o = wb_snoop[103];
  /* soc.vhdl:367:33  */
  assign n145_o = dmi_addr[3:0];
  /* soc.vhdl:269:26  */
  assign n154_o = n95_o[29:1];
  /* soc.vhdl:270:23  */
  assign n157_o = n95_o[61:30];
  /* soc.vhdl:270:32  */
  assign n158_o = n95_o[61:30];
  /* soc.vhdl:270:27  */
  assign n159_o = {n157_o, n158_o};
  /* soc.vhdl:272:18  */
  assign n163_o = n95_o[0];
  /* soc.vhdl:272:22  */
  assign n164_o = ~n163_o;
  /* soc.vhdl:273:39  */
  assign n165_o = n95_o[65:62];
  /* soc.vhdl:275:39  */
  assign n166_o = n95_o[65:62];
  assign n167_o = n161_o[3:0];
  /* soc.vhdl:272:9  */
  assign n168_o = n164_o ? n165_o : n167_o;
  assign n169_o = n161_o[7:4];
  /* soc.vhdl:272:9  */
  assign n170_o = n164_o ? n169_o : n166_o;
  /* soc.vhdl:277:23  */
  assign n172_o = n95_o[66];
  /* soc.vhdl:278:23  */
  assign n174_o = n95_o[67];
  /* soc.vhdl:279:22  */
  assign n176_o = n95_o[68];
  assign n177_o = {n176_o, n174_o, n172_o, n170_o, n168_o, n159_o, n154_o};
  assign n178_o = {wishbone_dcore_out, wishbone_icore_out, n177_o, wishbone_debug_out};
  /* soc.vhdl:381:39  */
  assign n179_o = wb_masters_in[263:198];
  /* soc.vhdl:382:39  */
  assign n180_o = wb_masters_in[197:132];
  /* soc.vhdl:383:60  */
  assign n182_o = wb_masters_in[131:66];
  /* soc.vhdl:383:82  */
  assign n183_o = n95_o[29:0];
  /* soc.vhdl:287:25  */
  assign n189_o = n182_o[64];
  /* soc.vhdl:288:27  */
  assign n193_o = n182_o[65];
  /* soc.vhdl:289:15  */
  assign n194_o = n183_o[0];
  /* soc.vhdl:289:19  */
  assign n195_o = ~n194_o;
  /* soc.vhdl:290:32  */
  assign n196_o = n182_o[31:0];
  /* soc.vhdl:292:32  */
  assign n197_o = n182_o[63:32];
  /* soc.vhdl:289:9  */
  assign n198_o = n195_o ? n196_o : n197_o;
  assign n199_o = {n193_o, n189_o, n198_o};
  /* soc.vhdl:384:39  */
  assign n200_o = wb_masters_in[65:0];
  /* soc.vhdl:385:5  */
  wishbone_arbiter_4 wishbone_arbiter_0 (
    .clk(system_clk),
    .rst(rst_wbar),
    .wb_masters_in(wb_masters_out),
    .wb_slave_in_dat(n204_o),
    .wb_slave_in_ack(n205_o),
    .wb_slave_in_stall(n206_o),
    .wb_masters_out(wishbone_arbiter_0_wb_masters_out),
    .wb_slave_out_adr(wishbone_arbiter_0_wb_slave_out_adr),
    .wb_slave_out_dat(wishbone_arbiter_0_wb_slave_out_dat),
    .wb_slave_out_sel(wishbone_arbiter_0_wb_slave_out_sel),
    .wb_slave_out_cyc(wishbone_arbiter_0_wb_slave_out_cyc),
    .wb_slave_out_stb(wishbone_arbiter_0_wb_slave_out_stb),
    .wb_slave_out_we(wishbone_arbiter_0_wb_slave_out_we));
  assign n202_o = {wishbone_arbiter_0_wb_slave_out_we, wishbone_arbiter_0_wb_slave_out_stb, wishbone_arbiter_0_wb_slave_out_cyc, wishbone_arbiter_0_wb_slave_out_sel, wishbone_arbiter_0_wb_slave_out_dat, wishbone_arbiter_0_wb_slave_out_adr};
  assign n204_o = wb_master_in[63:0];
  assign n205_o = wb_master_in[64];
  assign n206_o = wb_master_in[65];
  /* soc.vhdl:405:25  */
  assign n209_o = wb_master_in[65];
  assign n211_o = wb_master_out[102];
  /* soc.vhdl:405:9  */
  assign n212_o = n209_o ? 1'b0 : n211_o;
  assign n213_o = wb_master_out[103];
  assign n214_o = wb_master_out[101:0];
  /* soc.vhdl:427:40  */
  assign n219_o = wb_master_out[28:26];
  /* soc.vhdl:427:55  */
  assign n220_o = {n219_o, dram_at_0};
  /* soc.vhdl:429:15  */
  assign n223_o = n220_o & 4'b1111;
  /* soc.vhdl:429:15  */
  assign n224_o = n223_o == 4'b0000;
  /* soc.vhdl:431:15  */
  assign n227_o = n220_o & 4'b1111;
  /* soc.vhdl:431:15  */
  assign n228_o = n227_o == 4'b0001;
  /* soc.vhdl:433:15  */
  assign n231_o = n220_o & 4'b1100;
  /* soc.vhdl:433:15  */
  assign n232_o = n231_o == 4'b0100;
  /* soc.vhdl:435:15  */
  assign n235_o = n220_o & 4'b1100;
  /* soc.vhdl:435:15  */
  assign n236_o = n235_o == 4'b1000;
  /* soc.vhdl:437:15  */
  assign n239_o = n220_o & 4'b1100;
  /* soc.vhdl:437:15  */
  assign n240_o = n239_o == 4'b1100;
  /* soc.vhdl:437:9  */
  assign n243_o = n240_o ? 2'b10 : 2'b00;
  /* soc.vhdl:435:9  */
  assign n245_o = n236_o ? 2'b00 : n243_o;
  /* soc.vhdl:433:9  */
  assign n247_o = n232_o ? 2'b01 : n245_o;
  /* soc.vhdl:431:9  */
  assign n249_o = n228_o ? 2'b01 : n247_o;
  /* soc.vhdl:429:9  */
  assign n251_o = n224_o ? 2'b00 : n249_o;
  assign n254_o = wb_master_out[103:102];
  assign n255_o = wb_master_out[100:0];
  assign n257_o = wb_master_out[103:102];
  assign n258_o = wb_master_out[100:0];
  assign n260_o = wb_master_out[103:102];
  assign n261_o = wb_master_out[100:0];
  /* soc.vhdl:450:45  */
  assign n262_o = wb_master_out[101];
  /* soc.vhdl:449:9  */
  assign n264_o = n251_o == 2'b00;
  /* soc.vhdl:454:49  */
  assign n265_o = wb_master_out[101];
  /* soc.vhdl:452:9  */
  assign n267_o = n251_o == 2'b01;
  /* soc.vhdl:462:43  */
  assign n268_o = wb_master_out[101];
  /* soc.vhdl:461:9  */
  assign n270_o = n251_o == 2'b10;
  assign n271_o = {n270_o, n267_o, n264_o};
  /* soc.vhdl:448:9  */
  always @*
    case (n271_o)
      3'b100: n273_o = 1'b0;
      3'b010: n273_o = n265_o;
      3'b001: n273_o = 1'b0;
      default: n273_o = 1'bX;
    endcase
  /* soc.vhdl:448:9  */
  always @*
    case (n271_o)
      3'b100: n275_o = wb_io_out;
      3'b010: n275_o = n77_o;
      3'b001: n275_o = wb_bram_out;
      default: n275_o = 66'bX;
    endcase
  /* soc.vhdl:448:9  */
  always @*
    case (n271_o)
      3'b100: n277_o = n268_o;
      3'b010: n277_o = 1'b0;
      3'b001: n277_o = 1'b0;
      default: n277_o = 1'bX;
    endcase
  /* soc.vhdl:448:9  */
  always @*
    case (n271_o)
      3'b100: n279_o = 1'b0;
      3'b010: n279_o = 1'b0;
      3'b001: n279_o = n262_o;
      default: n279_o = 1'bX;
    endcase
  /* soc.vhdl:480:18  */
  always @*
    slave_io_latch_state = n756_q; // (isignal)
  initial
    slave_io_latch_state = 2'b00;
  /* soc.vhdl:483:18  */
  always @*
    slave_io_latch_has_top = n757_q; // (isignal)
  initial
    slave_io_latch_has_top = 1'b0;
  /* soc.vhdl:508:33  */
  assign n294_o = wb_io_in[101];
  /* soc.vhdl:508:56  */
  assign n295_o = wb_io_in[102];
  /* soc.vhdl:508:43  */
  assign n296_o = n294_o & n295_o;
  /* soc.vhdl:518:51  */
  assign n299_o = wb_io_in[103];
  /* soc.vhdl:519:55  */
  assign n300_o = wb_io_in[28:0];
  /* soc.vhdl:519:90  */
  assign n302_o = {n300_o, 1'b0};
  /* soc.vhdl:522:48  */
  assign n303_o = wb_io_in[100:97];
  /* soc.vhdl:522:61  */
  assign n305_o = n303_o != 4'b0000;
  /* soc.vhdl:523:48  */
  assign n306_o = wb_io_in[96:93];
  /* soc.vhdl:523:61  */
  assign n308_o = n306_o != 4'b0000;
  /* soc.vhdl:529:41  */
  assign n309_o = wb_io_in[103];
  /* soc.vhdl:530:63  */
  assign n310_o = wb_io_in[60:29];
  assign n311_o = wb_sio_out[61:30];
  /* soc.vhdl:529:29  */
  assign n312_o = n309_o ? n310_o : n311_o;
  /* soc.vhdl:532:59  */
  assign n313_o = wb_io_in[96:93];
  /* soc.vhdl:537:41  */
  assign n314_o = wb_io_in[103];
  /* soc.vhdl:538:63  */
  assign n315_o = wb_io_in[92:61];
  assign n316_o = wb_sio_out[61:30];
  /* soc.vhdl:537:29  */
  assign n317_o = n314_o ? n315_o : n316_o;
  /* soc.vhdl:540:59  */
  assign n318_o = wb_io_in[100:97];
  assign n320_o = {n318_o, n317_o};
  assign n321_o = {n313_o, n312_o};
  assign n322_o = n302_o[0];
  /* soc.vhdl:528:25  */
  assign n323_o = n308_o ? n322_o : 1'b1;
  /* soc.vhdl:528:25  */
  assign n324_o = n308_o ? n321_o : n320_o;
  assign n325_o = n302_o[29:1];
  /* soc.vhdl:528:25  */
  assign n328_o = n308_o ? 2'b01 : 2'b10;
  assign n329_o = wb_io_out[65];
  /* soc.vhdl:508:21  */
  assign n330_o = n296_o ? 1'b1 : n329_o;
  assign n331_o = {n324_o, n325_o, n323_o};
  assign n332_o = {n299_o, 1'b1};
  assign n333_o = wb_sio_out[65:0];
  /* soc.vhdl:508:21  */
  assign n334_o = n296_o ? n331_o : n333_o;
  assign n335_o = wb_sio_out[68:67];
  /* soc.vhdl:508:21  */
  assign n336_o = n296_o ? n332_o : n335_o;
  /* soc.vhdl:508:21  */
  assign n337_o = n296_o ? n328_o : slave_io_latch_state;
  /* soc.vhdl:508:21  */
  assign n338_o = n296_o ? n305_o : slave_io_latch_has_top;
  /* soc.vhdl:508:21  */
  assign n342_o = n296_o ? 1'b1 : 1'b0;
  /* soc.vhdl:503:17  */
  assign n344_o = slave_io_latch_state == 2'b00;
  /* soc.vhdl:551:34  */
  assign n345_o = wb_sio_in[33];
  /* soc.vhdl:551:40  */
  assign n346_o = ~n345_o;
  assign n348_o = wb_sio_out[67];
  /* soc.vhdl:551:21  */
  assign n349_o = n346_o ? 1'b0 : n348_o;
  /* soc.vhdl:556:34  */
  assign n350_o = wb_sio_in[32];
  /* soc.vhdl:558:39  */
  assign n351_o = wb_sio_out[68];
  /* soc.vhdl:558:42  */
  assign n352_o = ~n351_o;
  /* soc.vhdl:559:69  */
  assign n353_o = wb_sio_in[31:0];
  assign n354_o = wb_io_out[31:0];
  /* soc.vhdl:556:21  */
  assign n355_o = n381_o ? n353_o : n354_o;
  /* soc.vhdl:565:41  */
  assign n356_o = wb_io_in[103];
  /* soc.vhdl:566:63  */
  assign n357_o = wb_io_in[92:61];
  assign n358_o = wb_sio_out[61:30];
  /* soc.vhdl:565:29  */
  assign n359_o = n356_o ? n357_o : n358_o;
  /* soc.vhdl:568:59  */
  assign n360_o = wb_io_in[100:97];
  assign n365_o = {1'b0, 1'b1};
  assign n366_o = wb_io_out[65:64];
  /* soc.vhdl:563:25  */
  assign n367_o = slave_io_latch_has_top ? n366_o : n365_o;
  assign n368_o = {n360_o, n359_o};
  assign n369_o = wb_sio_out[0];
  /* soc.vhdl:556:21  */
  assign n370_o = n385_o ? 1'b1 : n369_o;
  assign n371_o = wb_sio_out[65:30];
  /* soc.vhdl:556:21  */
  assign n372_o = n387_o ? n368_o : n371_o;
  /* soc.vhdl:556:21  */
  assign n373_o = n388_o ? 1'b1 : n349_o;
  /* soc.vhdl:563:25  */
  assign n376_o = slave_io_latch_has_top ? 2'b10 : 2'b00;
  /* soc.vhdl:563:25  */
  assign n379_o = slave_io_latch_has_top ? 1'b0 : 1'b1;
  /* soc.vhdl:556:21  */
  assign n381_o = n350_o & n352_o;
  assign n382_o = wb_io_out[65:64];
  /* soc.vhdl:556:21  */
  assign n383_o = n350_o ? n367_o : n382_o;
  /* soc.vhdl:556:21  */
  assign n385_o = n350_o & slave_io_latch_has_top;
  /* soc.vhdl:556:21  */
  assign n387_o = n350_o & slave_io_latch_has_top;
  /* soc.vhdl:556:21  */
  assign n388_o = n350_o & slave_io_latch_has_top;
  /* soc.vhdl:556:21  */
  assign n389_o = n350_o ? n376_o : slave_io_latch_state;
  /* soc.vhdl:556:21  */
  assign n391_o = n350_o ? n379_o : 1'b0;
  /* soc.vhdl:549:17  */
  assign n393_o = slave_io_latch_state == 2'b01;
  /* soc.vhdl:590:34  */
  assign n394_o = wb_sio_in[33];
  /* soc.vhdl:590:40  */
  assign n395_o = ~n394_o;
  assign n397_o = wb_sio_out[67];
  /* soc.vhdl:590:21  */
  assign n398_o = n395_o ? 1'b0 : n397_o;
  /* soc.vhdl:595:34  */
  assign n399_o = wb_sio_in[32];
  /* soc.vhdl:597:39  */
  assign n400_o = wb_sio_out[68];
  /* soc.vhdl:597:42  */
  assign n401_o = ~n400_o;
  /* soc.vhdl:598:70  */
  assign n402_o = wb_sio_in[31:0];
  assign n403_o = wb_io_out[63:32];
  /* soc.vhdl:597:25  */
  assign n404_o = n401_o ? n402_o : n403_o;
  assign n407_o = {1'b0, 1'b1, n404_o};
  assign n408_o = wb_io_out[65:32];
  /* soc.vhdl:595:21  */
  assign n409_o = n399_o ? n407_o : n408_o;
  /* soc.vhdl:595:21  */
  assign n411_o = n399_o ? 2'b00 : slave_io_latch_state;
  /* soc.vhdl:595:21  */
  assign n414_o = n399_o ? 1'b1 : 1'b0;
  /* soc.vhdl:588:17  */
  assign n416_o = slave_io_latch_state == 2'b10;
  assign n417_o = {n416_o, n393_o, n344_o};
  assign n418_o = wb_io_out[31:0];
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n420_o = n418_o;
      3'b010: n420_o = n355_o;
      3'b001: n420_o = n418_o;
      default: n420_o = 32'bX;
    endcase
  assign n421_o = n409_o[31:0];
  assign n422_o = wb_io_out[63:32];
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n424_o = n421_o;
      3'b010: n424_o = n422_o;
      3'b001: n424_o = n422_o;
      default: n424_o = 32'bX;
    endcase
  assign n425_o = n383_o[0];
  assign n426_o = n409_o[32];
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n428_o = n426_o;
      3'b010: n428_o = n425_o;
      3'b001: n428_o = 1'b0;
      default: n428_o = 1'bX;
    endcase
  assign n429_o = n383_o[1];
  assign n430_o = n409_o[33];
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n432_o = n430_o;
      3'b010: n432_o = n429_o;
      3'b001: n432_o = n330_o;
      default: n432_o = 1'bX;
    endcase
  assign n433_o = n334_o[0];
  assign n434_o = wb_sio_out[0];
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n436_o = n434_o;
      3'b010: n436_o = n370_o;
      3'b001: n436_o = n433_o;
      default: n436_o = 1'bX;
    endcase
  assign n437_o = n334_o[29:1];
  assign n438_o = wb_sio_out[29:1];
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n440_o = n438_o;
      3'b010: n440_o = n438_o;
      3'b001: n440_o = n437_o;
      default: n440_o = 29'bX;
    endcase
  assign n441_o = n334_o[65:30];
  assign n442_o = wb_sio_out[65:30];
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n444_o = n442_o;
      3'b010: n444_o = n372_o;
      3'b001: n444_o = n441_o;
      default: n444_o = 36'bX;
    endcase
  assign n445_o = n336_o[0];
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n447_o = n398_o;
      3'b010: n447_o = n373_o;
      3'b001: n447_o = n445_o;
      default: n447_o = 1'bX;
    endcase
  assign n448_o = n336_o[1];
  assign n449_o = wb_sio_out[68];
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n451_o = n449_o;
      3'b010: n451_o = n449_o;
      3'b001: n451_o = n448_o;
      default: n451_o = 1'bX;
    endcase
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n453_o = n411_o;
      3'b010: n453_o = n389_o;
      3'b001: n453_o = n337_o;
      default: n453_o = 2'bX;
    endcase
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n455_o = slave_io_latch_has_top;
      3'b010: n455_o = slave_io_latch_has_top;
      3'b001: n455_o = n338_o;
      default: n455_o = 1'bX;
    endcase
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n460_o = 1'b0;
      3'b010: n460_o = 1'b0;
      3'b001: n460_o = n342_o;
      default: n460_o = 1'bX;
    endcase
  /* soc.vhdl:502:17  */
  always @*
    case (n417_o)
      3'b100: n463_o = n414_o;
      3'b010: n463_o = n391_o;
      3'b001: n463_o = 1'b0;
      default: n463_o = 1'bX;
    endcase
  assign n464_o = {n432_o, n428_o, n424_o, n420_o};
  assign n465_o = {1'b0, 1'b0};
  assign n466_o = n464_o[63:0];
  assign n467_o = wb_io_out[63:0];
  /* soc.vhdl:493:13  */
  assign n468_o = rst ? n467_o : n466_o;
  assign n469_o = n464_o[65:64];
  /* soc.vhdl:493:13  */
  assign n470_o = rst ? n465_o : n469_o;
  assign n471_o = {n444_o, n440_o, n436_o};
  assign n472_o = {n451_o, n447_o};
  assign n473_o = wb_sio_out[65:0];
  /* soc.vhdl:493:13  */
  assign n474_o = rst ? n473_o : n471_o;
  assign n475_o = n472_o[0];
  /* soc.vhdl:493:13  */
  assign n476_o = rst ? 1'b0 : n475_o;
  assign n477_o = n472_o[1];
  assign n478_o = wb_sio_out[68];
  /* soc.vhdl:493:13  */
  assign n479_o = rst ? n478_o : n477_o;
  /* soc.vhdl:493:13  */
  assign n481_o = rst ? 2'b00 : n453_o;
  /* soc.vhdl:493:13  */
  assign n483_o = rst ? 1'b0 : n455_o;
  /* soc.vhdl:493:13  */
  assign n487_o = rst ? 1'b0 : n460_o;
  /* soc.vhdl:493:13  */
  assign n490_o = rst ? 1'b1 : n463_o;
  /* soc.vhdl:616:29  */
  assign n492_o = n487_o | n490_o;
  /* soc.vhdl:616:13  */
  assign n495_o = n492_o ? 1'b0 : n997_q;
  /* soc.vhdl:616:13  */
  assign n497_o = n492_o ? 1'b0 : n998_q;
  assign n502_o = wb_sio_out[66];
  /* soc.vhdl:616:13  */
  assign n503_o = n492_o ? 1'b0 : n502_o;
  /* soc.vhdl:616:13  */
  assign n505_o = n492_o ? 1'b0 : wb_spiflash_is_reg;
  /* soc.vhdl:616:13  */
  assign n507_o = n492_o ? 1'b0 : wb_spiflash_is_map;
  /* soc.vhdl:616:13  */
  assign n509_o = n492_o ? 1'b0 : io_cycle_none;
  /* soc.vhdl:616:13  */
  assign n511_o = n492_o ? 1'b0 : io_cycle_syscon;
  /* soc.vhdl:616:13  */
  assign n513_o = n492_o ? 1'b0 : io_cycle_uart;
  /* soc.vhdl:616:13  */
  assign n515_o = n492_o ? 1'b0 : io_cycle_uart1;
  /* soc.vhdl:616:13  */
  assign n517_o = n492_o ? 1'b0 : io_cycle_icp;
  /* soc.vhdl:616:13  */
  assign n519_o = n492_o ? 1'b0 : io_cycle_ics;
  /* soc.vhdl:616:13  */
  assign n521_o = n492_o ? 1'b0 : io_cycle_spi_flash;
  /* soc.vhdl:616:13  */
  assign n523_o = n492_o ? 1'b0 : io_cycle_gpio;
  /* soc.vhdl:616:13  */
  assign n525_o = n492_o ? 1'b0 : io_cycle_external;
  /* soc.vhdl:637:45  */
  assign n526_o = wb_io_in[26:9];
  /* soc.vhdl:637:31  */
  assign n528_o = {2'b11, n526_o};
  /* soc.vhdl:639:23  */
  assign n531_o = n528_o & 20'b11111111000000000000;
  /* soc.vhdl:639:23  */
  assign n532_o = n531_o == 20'b11111111000000000000;
  /* soc.vhdl:639:50  */
  assign n534_o = n532_o & 1'b1;
  /* soc.vhdl:643:23  */
  assign n537_o = n528_o & 20'b11110000000000000000;
  /* soc.vhdl:643:23  */
  assign n538_o = n537_o == 20'b11110000000000000000;
  /* soc.vhdl:647:23  */
  assign n541_o = n528_o & 20'b11111111000000000000;
  /* soc.vhdl:647:23  */
  assign n542_o = n541_o == 20'b11001000000000000000;
  /* soc.vhdl:649:27  */
  assign n545_o = n528_o & 20'b00000000111111110000;
  /* soc.vhdl:649:27  */
  assign n546_o = n545_o == 20'b00000000000000000000;
  /* soc.vhdl:649:54  */
  assign n548_o = n546_o & 1'b1;
  /* soc.vhdl:647:17  */
  assign n563_o = n664_o ? 1'b1 : n495_o;
  /* soc.vhdl:649:21  */
  assign n565_o = n548_o ? n509_o : 1'b1;
  /* soc.vhdl:647:17  */
  assign n567_o = n674_o ? 1'b1 : n525_o;
  /* soc.vhdl:649:21  */
  assign n570_o = n548_o ? 3'b111 : 3'b000;
  /* soc.vhdl:665:23  */
  assign n573_o = n528_o & 20'b11111111111111111111;
  /* soc.vhdl:665:23  */
  assign n574_o = n573_o == 20'b11000000000000000000;
  /* soc.vhdl:668:23  */
  assign n577_o = n528_o & 20'b11111111111111111111;
  /* soc.vhdl:668:23  */
  assign n578_o = n577_o == 20'b11000000000000000010;
  /* soc.vhdl:671:23  */
  assign n581_o = n528_o & 20'b11111111111111111111;
  /* soc.vhdl:671:23  */
  assign n582_o = n581_o == 20'b11000000000000000011;
  /* soc.vhdl:674:23  */
  assign n585_o = n528_o & 20'b11111111111111111111;
  /* soc.vhdl:674:23  */
  assign n586_o = n585_o == 20'b11000000000000000100;
  /* soc.vhdl:677:23  */
  assign n589_o = n528_o & 20'b11111111111111111111;
  /* soc.vhdl:677:23  */
  assign n590_o = n589_o == 20'b11000000000000000101;
  /* soc.vhdl:680:23  */
  assign n593_o = n528_o & 20'b11111111111111111111;
  /* soc.vhdl:680:23  */
  assign n594_o = n593_o == 20'b11000000000000000110;
  /* soc.vhdl:684:23  */
  assign n597_o = n528_o & 20'b11111111111111111111;
  /* soc.vhdl:684:23  */
  assign n598_o = n597_o == 20'b11000000000000000111;
  /* soc.vhdl:684:17  */
  assign n600_o = n598_o ? n509_o : 1'b1;
  /* soc.vhdl:684:17  */
  assign n602_o = n598_o ? 1'b1 : n523_o;
  /* soc.vhdl:684:17  */
  assign n605_o = n598_o ? 3'b110 : 3'b000;
  /* soc.vhdl:680:17  */
  assign n607_o = n594_o ? 1'b1 : n505_o;
  /* soc.vhdl:680:17  */
  assign n608_o = n594_o ? n509_o : n600_o;
  /* soc.vhdl:680:17  */
  assign n610_o = n594_o ? 1'b1 : n521_o;
  /* soc.vhdl:680:17  */
  assign n611_o = n594_o ? n523_o : n602_o;
  /* soc.vhdl:680:17  */
  assign n613_o = n594_o ? 3'b101 : n605_o;
  /* soc.vhdl:677:17  */
  assign n614_o = n590_o ? n505_o : n607_o;
  /* soc.vhdl:677:17  */
  assign n615_o = n590_o ? n509_o : n608_o;
  /* soc.vhdl:677:17  */
  assign n617_o = n590_o ? 1'b1 : n519_o;
  /* soc.vhdl:677:17  */
  assign n618_o = n590_o ? n521_o : n610_o;
  /* soc.vhdl:677:17  */
  assign n619_o = n590_o ? n523_o : n611_o;
  /* soc.vhdl:677:17  */
  assign n621_o = n590_o ? 3'b011 : n613_o;
  /* soc.vhdl:674:17  */
  assign n622_o = n586_o ? n505_o : n614_o;
  /* soc.vhdl:674:17  */
  assign n623_o = n586_o ? n509_o : n615_o;
  /* soc.vhdl:674:17  */
  assign n625_o = n586_o ? 1'b1 : n517_o;
  /* soc.vhdl:674:17  */
  assign n626_o = n586_o ? n519_o : n617_o;
  /* soc.vhdl:674:17  */
  assign n627_o = n586_o ? n521_o : n618_o;
  /* soc.vhdl:674:17  */
  assign n628_o = n586_o ? n523_o : n619_o;
  /* soc.vhdl:674:17  */
  assign n630_o = n586_o ? 3'b010 : n621_o;
  /* soc.vhdl:671:17  */
  assign n631_o = n582_o ? n505_o : n622_o;
  /* soc.vhdl:671:17  */
  assign n632_o = n582_o ? n509_o : n623_o;
  /* soc.vhdl:671:17  */
  assign n634_o = n582_o ? 1'b1 : n515_o;
  /* soc.vhdl:671:17  */
  assign n635_o = n582_o ? n517_o : n625_o;
  /* soc.vhdl:671:17  */
  assign n636_o = n582_o ? n519_o : n626_o;
  /* soc.vhdl:671:17  */
  assign n637_o = n582_o ? n521_o : n627_o;
  /* soc.vhdl:671:17  */
  assign n638_o = n582_o ? n523_o : n628_o;
  /* soc.vhdl:671:17  */
  assign n640_o = n582_o ? 3'b100 : n630_o;
  /* soc.vhdl:668:17  */
  assign n641_o = n578_o ? n505_o : n631_o;
  /* soc.vhdl:668:17  */
  assign n642_o = n578_o ? n509_o : n632_o;
  /* soc.vhdl:668:17  */
  assign n644_o = n578_o ? 1'b1 : n513_o;
  /* soc.vhdl:668:17  */
  assign n645_o = n578_o ? n515_o : n634_o;
  /* soc.vhdl:668:17  */
  assign n646_o = n578_o ? n517_o : n635_o;
  /* soc.vhdl:668:17  */
  assign n647_o = n578_o ? n519_o : n636_o;
  /* soc.vhdl:668:17  */
  assign n648_o = n578_o ? n521_o : n637_o;
  /* soc.vhdl:668:17  */
  assign n649_o = n578_o ? n523_o : n638_o;
  /* soc.vhdl:668:17  */
  assign n651_o = n578_o ? 3'b001 : n640_o;
  /* soc.vhdl:665:17  */
  assign n652_o = n574_o ? n505_o : n641_o;
  /* soc.vhdl:665:17  */
  assign n653_o = n574_o ? n509_o : n642_o;
  /* soc.vhdl:665:17  */
  assign n655_o = n574_o ? 1'b1 : n511_o;
  /* soc.vhdl:665:17  */
  assign n656_o = n574_o ? n513_o : n644_o;
  /* soc.vhdl:665:17  */
  assign n657_o = n574_o ? n515_o : n645_o;
  /* soc.vhdl:665:17  */
  assign n658_o = n574_o ? n517_o : n646_o;
  /* soc.vhdl:665:17  */
  assign n659_o = n574_o ? n519_o : n647_o;
  /* soc.vhdl:665:17  */
  assign n660_o = n574_o ? n521_o : n648_o;
  /* soc.vhdl:665:17  */
  assign n661_o = n574_o ? n523_o : n649_o;
  /* soc.vhdl:665:17  */
  assign n663_o = n574_o ? 3'b000 : n651_o;
  /* soc.vhdl:647:17  */
  assign n664_o = n542_o & n548_o;
  /* soc.vhdl:647:17  */
  assign n665_o = n542_o ? n505_o : n652_o;
  /* soc.vhdl:647:17  */
  assign n666_o = n542_o ? n565_o : n653_o;
  /* soc.vhdl:647:17  */
  assign n667_o = n542_o ? n511_o : n655_o;
  /* soc.vhdl:647:17  */
  assign n668_o = n542_o ? n513_o : n656_o;
  /* soc.vhdl:647:17  */
  assign n669_o = n542_o ? n515_o : n657_o;
  /* soc.vhdl:647:17  */
  assign n670_o = n542_o ? n517_o : n658_o;
  /* soc.vhdl:647:17  */
  assign n671_o = n542_o ? n519_o : n659_o;
  /* soc.vhdl:647:17  */
  assign n672_o = n542_o ? n521_o : n660_o;
  /* soc.vhdl:647:17  */
  assign n673_o = n542_o ? n523_o : n661_o;
  /* soc.vhdl:647:17  */
  assign n674_o = n542_o & n548_o;
  /* soc.vhdl:647:17  */
  assign n675_o = n542_o ? n570_o : n663_o;
  /* soc.vhdl:643:17  */
  assign n676_o = n538_o ? n495_o : n563_o;
  /* soc.vhdl:643:17  */
  assign n677_o = n538_o ? n505_o : n665_o;
  /* soc.vhdl:643:17  */
  assign n679_o = n538_o ? 1'b1 : n507_o;
  /* soc.vhdl:643:17  */
  assign n680_o = n538_o ? n509_o : n666_o;
  /* soc.vhdl:643:17  */
  assign n681_o = n538_o ? n511_o : n667_o;
  /* soc.vhdl:643:17  */
  assign n682_o = n538_o ? n513_o : n668_o;
  /* soc.vhdl:643:17  */
  assign n683_o = n538_o ? n515_o : n669_o;
  /* soc.vhdl:643:17  */
  assign n684_o = n538_o ? n517_o : n670_o;
  /* soc.vhdl:643:17  */
  assign n685_o = n538_o ? n519_o : n671_o;
  /* soc.vhdl:643:17  */
  assign n687_o = n538_o ? 1'b1 : n672_o;
  /* soc.vhdl:643:17  */
  assign n688_o = n538_o ? n523_o : n673_o;
  /* soc.vhdl:643:17  */
  assign n689_o = n538_o ? n525_o : n567_o;
  /* soc.vhdl:643:17  */
  assign n691_o = n538_o ? 3'b101 : n675_o;
  /* soc.vhdl:639:17  */
  assign n692_o = n534_o ? n495_o : n676_o;
  /* soc.vhdl:634:13  */
  assign n694_o = n712_o ? 1'b1 : n497_o;
  /* soc.vhdl:639:17  */
  assign n695_o = n534_o ? n505_o : n677_o;
  /* soc.vhdl:639:17  */
  assign n696_o = n534_o ? n507_o : n679_o;
  /* soc.vhdl:639:17  */
  assign n697_o = n534_o ? n509_o : n680_o;
  /* soc.vhdl:639:17  */
  assign n698_o = n534_o ? n511_o : n681_o;
  /* soc.vhdl:639:17  */
  assign n699_o = n534_o ? n513_o : n682_o;
  /* soc.vhdl:639:17  */
  assign n700_o = n534_o ? n515_o : n683_o;
  /* soc.vhdl:639:17  */
  assign n701_o = n534_o ? n517_o : n684_o;
  /* soc.vhdl:639:17  */
  assign n702_o = n534_o ? n519_o : n685_o;
  /* soc.vhdl:639:17  */
  assign n703_o = n534_o ? n521_o : n687_o;
  /* soc.vhdl:639:17  */
  assign n704_o = n534_o ? n523_o : n688_o;
  /* soc.vhdl:639:17  */
  assign n706_o = n534_o ? 1'b1 : n689_o;
  /* soc.vhdl:639:17  */
  assign n708_o = n534_o ? 3'b111 : n691_o;
  /* soc.vhdl:634:13  */
  assign n711_o = n487_o ? n692_o : n495_o;
  /* soc.vhdl:634:13  */
  assign n712_o = n487_o & n534_o;
  /* soc.vhdl:634:13  */
  assign n713_o = n487_o ? 1'b1 : n503_o;
  /* soc.vhdl:634:13  */
  assign n714_o = n487_o ? n695_o : n505_o;
  /* soc.vhdl:634:13  */
  assign n715_o = n487_o ? n696_o : n507_o;
  /* soc.vhdl:634:13  */
  assign n717_o = n487_o ? n697_o : n509_o;
  /* soc.vhdl:634:13  */
  assign n718_o = n487_o ? n698_o : n511_o;
  /* soc.vhdl:634:13  */
  assign n719_o = n487_o ? n699_o : n513_o;
  /* soc.vhdl:634:13  */
  assign n720_o = n487_o ? n700_o : n515_o;
  /* soc.vhdl:634:13  */
  assign n721_o = n487_o ? n701_o : n517_o;
  /* soc.vhdl:634:13  */
  assign n722_o = n487_o ? n702_o : n519_o;
  /* soc.vhdl:634:13  */
  assign n723_o = n487_o ? n703_o : n521_o;
  /* soc.vhdl:634:13  */
  assign n724_o = n487_o ? n704_o : n523_o;
  /* soc.vhdl:634:13  */
  assign n725_o = n487_o ? n706_o : n525_o;
  assign n732_o = {n470_o, n468_o};
  assign n734_o = {n479_o, n476_o, n713_o, n474_o};
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n756_q <= n481_o;
  initial
    n756_q = 2'b00;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n757_q <= n483_o;
  initial
    n757_q = 1'b0;
  assign n760_o = wb_sio_out[68:67];
  assign n761_o = wb_sio_out[65:0];
  assign n762_o = wb_sio_out[68:67];
  assign n763_o = wb_sio_out[65:0];
  assign n764_o = wb_sio_out[68:67];
  assign n767_o = wb_sio_out[65:28];
  assign n768_o = wb_sio_out[25:0];
  assign n769_o = wb_sio_out[68:67];
  assign n770_o = wb_sio_out[65:0];
  /* soc.vhdl:717:57  */
  assign n773_o = wb_sio_out[5:0];
  assign n774_o = n771_o[29:6];
  assign n775_o = wb_sio_out[68:67];
  assign n776_o = wb_sio_out[65:30];
  /* soc.vhdl:721:57  */
  assign n779_o = wb_sio_out[9:0];
  assign n780_o = n777_o[29:10];
  assign n781_o = wb_sio_out[68:67];
  assign n782_o = wb_sio_out[65:30];
  assign n783_o = wb_sio_out[68:67];
  assign n784_o = wb_sio_out[65:0];
  assign n785_o = wb_sio_out[68:67];
  assign n786_o = wb_sio_out[65:0];
  /* soc.vhdl:731:9  */
  assign n788_o = current_io_decode == 3'b111;
  /* soc.vhdl:733:9  */
  assign n790_o = current_io_decode == 3'b000;
  /* soc.vhdl:735:9  */
  assign n792_o = current_io_decode == 3'b001;
  /* soc.vhdl:737:9  */
  assign n794_o = current_io_decode == 3'b010;
  /* soc.vhdl:739:9  */
  assign n796_o = current_io_decode == 3'b011;
  /* soc.vhdl:741:9  */
  assign n798_o = current_io_decode == 3'b100;
  /* soc.vhdl:743:9  */
  assign n800_o = current_io_decode == 3'b101;
  /* soc.vhdl:745:9  */
  assign n802_o = current_io_decode == 3'b110;
  assign n803_o = {n802_o, n800_o, n798_o, n796_o, n794_o, n792_o, n790_o, n788_o};
  /* soc.vhdl:730:9  */
  always @*
    case (n803_o)
      8'b10000000: n805_o = wb_gpio_out;
      8'b01000000: n805_o = wb_spiflash_out;
      8'b00100000: n805_o = wb_uart1_out;
      8'b00010000: n805_o = wb_xics_ics_out;
      8'b00001000: n805_o = wb_xics_icp_out;
      8'b00000100: n805_o = wb_uart0_out;
      8'b00000010: n805_o = wb_syscon_out;
      8'b00000001: n805_o = n85_o;
      default: n805_o = 34'bX;
    endcase
  /* soc.vhdl:752:41  */
  assign n807_o = wb_sio_out[67];
  /* soc.vhdl:752:60  */
  assign n808_o = wb_sio_out[66];
  /* soc.vhdl:752:45  */
  assign n809_o = n807_o & n808_o;
  assign n811_o = {1'b0, n809_o, 32'b11111111111111111111111111111111};
  /* soc.vhdl:750:9  */
  assign n812_o = io_cycle_none ? n811_o : n805_o;
  /* soc.vhdl:759:5  */
  syscon_100000000_4096_0_0_0_589433b711fb88bdee7cbb7d486960b51e4c8efd syscon0 (
    .clk(system_clk),
    .rst(rst),
    .wishbone_in_adr(n814_o),
    .wishbone_in_dat(n815_o),
    .wishbone_in_sel(n816_o),
    .wishbone_in_cyc(n817_o),
    .wishbone_in_stb(n818_o),
    .wishbone_in_we(n819_o),
    .wishbone_out_dat(syscon0_wishbone_out_dat),
    .wishbone_out_ack(syscon0_wishbone_out_ack),
    .wishbone_out_stall(syscon0_wishbone_out_stall),
    .dram_at_0(syscon0_dram_at_0),
    .core_reset(syscon0_core_reset),
    .soc_reset());
  assign n814_o = wb_syscon_in[29:0];
  assign n815_o = wb_syscon_in[61:30];
  assign n816_o = wb_syscon_in[65:62];
  assign n817_o = wb_syscon_in[66];
  assign n818_o = wb_syscon_in[67];
  assign n819_o = wb_syscon_in[68];
  assign n820_o = {syscon0_wishbone_out_stall, syscon0_wishbone_out_ack, syscon0_wishbone_out_dat};
  /* soc.vhdl:811:16  */
  assign uart0_16550_irq_l = uart0_16550_uart0_int_o; // (signal)
  /* soc.vhdl:813:9  */
  uart_top uart0_16550_uart0 (
    .wb_clk_i(system_clk),
    .wb_rst_i(rst_uart),
    .wb_adr_i(n824_o),
    .wb_dat_i(n825_o),
    .wb_we_i(n827_o),
    .wb_stb_i(n828_o),
    .wb_cyc_i(n829_o),
    .srx_pad_i(uart0_rxd),
    .cts_pad_i(n833_o),
    .dsr_pad_i(n834_o),
    .ri_pad_i(n835_o),
    .dcd_pad_i(n836_o),
    .wb_dat_o(uart0_16550_uart0_wb_dat_o),
    .wb_ack_o(uart0_16550_uart0_wb_ack_o),
    .int_o(uart0_16550_uart0_int_o),
    .stx_pad_o(uart0_16550_uart0_stx_pad_o),
    .rts_pad_o(),
    .dtr_pad_o());
  /* soc.vhdl:817:46  */
  assign n824_o = wb_uart0_in[2:0];
  /* soc.vhdl:818:46  */
  assign n825_o = wb_uart0_in[37:30];
  /* soc.vhdl:820:43  */
  assign n827_o = wb_uart0_in[68];
  /* soc.vhdl:821:43  */
  assign n828_o = wb_uart0_in[67];
  /* soc.vhdl:822:43  */
  assign n829_o = wb_uart0_in[66];
  /* soc.vhdl:844:35  */
  assign n842_o = {24'b000000000000000000000000, uart0_dat8};
  /* soc.vhdl:845:44  */
  assign n843_o = wb_uart0_out[32];
  /* soc.vhdl:845:27  */
  assign n844_o = ~n843_o;
  /* soc.vhdl:889:41  */
  assign n846_o = wb_uart1_in[66];
  /* soc.vhdl:889:61  */
  assign n847_o = wb_uart1_in[67];
  /* soc.vhdl:889:45  */
  assign n848_o = n846_o & n847_o;
  /* soc.vhdl:895:9  */
  spi_flash_ctrl_4_4_1489f923c4dca729178b3e3233458550d8dddf29 spiflash_gen_spiflash (
    .clk(system_clk),
    .rst(rst_spi),
    .wb_in_adr(n851_o),
    .wb_in_dat(n852_o),
    .wb_in_sel(n853_o),
    .wb_in_cyc(n854_o),
    .wb_in_stb(n855_o),
    .wb_in_we(n856_o),
    .wb_sel_reg(wb_spiflash_is_reg),
    .wb_sel_map(wb_spiflash_is_map),
    .sdat_i(spi_flash_sdat_i),
    .wb_out_dat(spiflash_gen_spiflash_wb_out_dat),
    .wb_out_ack(spiflash_gen_spiflash_wb_out_ack),
    .wb_out_stall(spiflash_gen_spiflash_wb_out_stall),
    .sck(spiflash_gen_spiflash_sck),
    .cs_n(spiflash_gen_spiflash_cs_n),
    .sdat_o(spiflash_gen_spiflash_sdat_o),
    .sdat_oe(spiflash_gen_spiflash_sdat_oe));
  assign n851_o = wb_spiflash_in[29:0];
  assign n852_o = wb_spiflash_in[61:30];
  assign n853_o = wb_spiflash_in[65:62];
  assign n854_o = wb_spiflash_in[66];
  assign n855_o = wb_spiflash_in[67];
  assign n856_o = wb_spiflash_in[68];
  assign n857_o = {spiflash_gen_spiflash_wb_out_stall, spiflash_gen_spiflash_wb_out_ack, spiflash_gen_spiflash_wb_out_dat};
  /* soc.vhdl:923:5  */
  xics_icp xics_icp (
    .clk(system_clk),
    .rst(rst_xics),
    .wb_in_adr(n863_o),
    .wb_in_dat(n864_o),
    .wb_in_sel(n865_o),
    .wb_in_cyc(n866_o),
    .wb_in_stb(n867_o),
    .wb_in_we(n868_o),
    .ics_in_src(n871_o),
    .ics_in_pri(n872_o),
    .wb_out_dat(xics_icp_wb_out_dat),
    .wb_out_ack(xics_icp_wb_out_ack),
    .wb_out_stall(xics_icp_wb_out_stall),
    .core_irq_out(xics_icp_core_irq_out));
  assign n863_o = wb_xics_icp_in[29:0];
  assign n864_o = wb_xics_icp_in[61:30];
  assign n865_o = wb_xics_icp_in[65:62];
  assign n866_o = wb_xics_icp_in[66];
  assign n867_o = wb_xics_icp_in[67];
  assign n868_o = wb_xics_icp_in[68];
  assign n869_o = {xics_icp_wb_out_stall, xics_icp_wb_out_ack, xics_icp_wb_out_dat};
  assign n871_o = ics_to_icp[3:0];
  assign n872_o = ics_to_icp[11:4];
  /* soc.vhdl:933:5  */
  xics_ics_16_3 xics_ics (
    .clk(system_clk),
    .rst(rst_xics),
    .wb_in_adr(n874_o),
    .wb_in_dat(n875_o),
    .wb_in_sel(n876_o),
    .wb_in_cyc(n877_o),
    .wb_in_stb(n878_o),
    .wb_in_we(n879_o),
    .int_level_in(int_level_in),
    .wb_out_dat(xics_ics_wb_out_dat),
    .wb_out_ack(xics_ics_wb_out_ack),
    .wb_out_stall(xics_ics_wb_out_stall),
    .icp_out_src(xics_ics_icp_out_src),
    .icp_out_pri(xics_ics_icp_out_pri));
  assign n874_o = wb_xics_ics_in[29:0];
  assign n875_o = wb_xics_ics_in[61:30];
  assign n876_o = wb_xics_ics_in[65:62];
  assign n877_o = wb_xics_ics_in[66];
  assign n878_o = wb_xics_ics_in[67];
  assign n879_o = wb_xics_ics_in[68];
  assign n880_o = {xics_ics_wb_out_stall, xics_ics_wb_out_ack, xics_ics_wb_out_dat};
  assign n882_o = {xics_ics_icp_out_pri, xics_ics_icp_out_src};
  /* soc.vhdl:948:9  */
  gpio_32 gpio0_gen_gpio (
    .clk(system_clk),
    .rst(rst_gpio),
    .wb_in_adr(n884_o),
    .wb_in_dat(n885_o),
    .wb_in_sel(n886_o),
    .wb_in_cyc(n887_o),
    .wb_in_stb(n888_o),
    .wb_in_we(n889_o),
    .gpio_in(gpio_in),
    .wb_out_dat(gpio0_gen_gpio_wb_out_dat),
    .wb_out_ack(gpio0_gen_gpio_wb_out_ack),
    .wb_out_stall(gpio0_gen_gpio_wb_out_stall),
    .gpio_out(gpio0_gen_gpio_gpio_out),
    .gpio_dir(gpio0_gen_gpio_gpio_dir),
    .intr(gpio0_gen_gpio_intr));
  assign n884_o = wb_gpio_in[29:0];
  assign n885_o = wb_gpio_in[61:30];
  assign n886_o = wb_gpio_in[65:62];
  assign n887_o = wb_gpio_in[66];
  assign n888_o = wb_gpio_in[67];
  assign n889_o = wb_gpio_in[68];
  assign n890_o = {gpio0_gen_gpio_wb_out_stall, gpio0_gen_gpio_wb_out_ack, gpio0_gen_gpio_wb_out_dat};
  assign n901_o = n896_o[15:5];
  /* soc.vhdl:977:9  */
  wishbone_bram_wrapper_4096_a75adb9e07879fb6c63b494abe06e3f9a6bb2ed9 bram_bram0 (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .clk(system_clk),
    .rst(rst_bram),
    .wishbone_in_adr(n903_o),
    .wishbone_in_dat(n904_o),
    .wishbone_in_sel(n905_o),
    .wishbone_in_cyc(n906_o),
    .wishbone_in_stb(n907_o),
    .wishbone_in_we(n908_o),
    .wishbone_out_dat(bram_bram0_wishbone_out_dat),
    .wishbone_out_ack(bram_bram0_wishbone_out_ack),
    .wishbone_out_stall(bram_bram0_wishbone_out_stall));
  assign n903_o = wb_bram_in[28:0];
  assign n904_o = wb_bram_in[92:29];
  assign n905_o = wb_bram_in[100:93];
  assign n906_o = wb_bram_in[101];
  assign n907_o = wb_bram_in[102];
  assign n908_o = wb_bram_in[103];
  assign n909_o = {bram_bram0_wishbone_out_stall, bram_bram0_wishbone_out_ack, bram_bram0_wishbone_out_dat};
  /* soc.vhdl:998:9  */
  dmi_dtm_jtag_8_64 dmi_jtag_dtm (
    .sys_clk(system_clk),
    .sys_reset(rst_dtm),
    .dmi_din(dmi_din),
    .dmi_ack(dmi_ack),
    .jtag_tck(jtag_tck),
    .jtag_tdi(jtag_tdi),
    .jtag_tms(jtag_tms),
    .jtag_trst(jtag_trst),
    .dmi_addr(dmi_jtag_dtm_dmi_addr),
    .dmi_dout(dmi_jtag_dtm_dmi_dout),
    .dmi_req(dmi_jtag_dtm_dmi_req),
    .dmi_wr(dmi_jtag_dtm_dmi_wr),
    .jtag_tdo(dmi_jtag_dtm_jtag_tdo));
  /* soc.vhdl:1056:12  */
  assign n920_o = dmi_addr & 8'b11111100;
  /* soc.vhdl:1056:12  */
  assign n921_o = n920_o == 8'b00000000;
  /* soc.vhdl:1058:15  */
  assign n924_o = dmi_addr & 8'b11110000;
  /* soc.vhdl:1058:15  */
  assign n925_o = n924_o == 8'b00010000;
  /* soc.vhdl:1058:9  */
  assign n928_o = n925_o ? 2'b01 : 2'b10;
  /* soc.vhdl:1056:9  */
  assign n930_o = n921_o ? 2'b00 : n928_o;
  /* soc.vhdl:1066:9  */
  assign n933_o = n930_o == 2'b00;
  /* soc.vhdl:1070:9  */
  assign n935_o = n930_o == 2'b01;
  assign n936_o = {n935_o, n933_o};
  /* soc.vhdl:1065:9  */
  always @*
    case (n936_o)
      2'b10: n938_o = dmi_core_dout;
      2'b01: n938_o = dmi_wb_dout;
      default: n938_o = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    endcase
  /* soc.vhdl:1065:9  */
  always @*
    case (n936_o)
      2'b10: n939_o = dmi_core_ack;
      2'b01: n939_o = dmi_wb_ack;
      default: n939_o = dmi_req;
    endcase
  /* soc.vhdl:1065:9  */
  always @*
    case (n936_o)
      2'b10: n941_o = 1'b0;
      2'b01: n941_o = dmi_req;
      default: n941_o = 1'b0;
    endcase
  /* soc.vhdl:1065:9  */
  always @*
    case (n936_o)
      2'b10: n944_o = dmi_req;
      2'b01: n944_o = 1'b0;
      default: n944_o = 1'b0;
    endcase
  /* soc.vhdl:1086:5  */
  wishbone_debug_master wishbone_debug (
    .clk(system_clk),
    .rst(rst_wbdb),
    .dmi_addr(n947_o),
    .dmi_din(dmi_dout),
    .dmi_req(dmi_wb_req),
    .dmi_wr(dmi_wr),
    .wb_in_dat(n952_o),
    .wb_in_ack(n953_o),
    .wb_in_stall(n954_o),
    .dmi_dout(wishbone_debug_dmi_dout),
    .dmi_ack(wishbone_debug_dmi_ack),
    .wb_out_adr(wishbone_debug_wb_out_adr),
    .wb_out_dat(wishbone_debug_wb_out_dat),
    .wb_out_sel(wishbone_debug_wb_out_sel),
    .wb_out_cyc(wishbone_debug_wb_out_cyc),
    .wb_out_stb(wishbone_debug_wb_out_stb),
    .wb_out_we(wishbone_debug_wb_out_we));
  /* soc.vhdl:1089:38  */
  assign n947_o = dmi_addr[1:0];
  assign n950_o = {wishbone_debug_wb_out_we, wishbone_debug_wb_out_stb, wishbone_debug_wb_out_cyc, wishbone_debug_wb_out_sel, wishbone_debug_wb_out_dat, wishbone_debug_wb_out_adr};
  assign n952_o = wishbone_debug_in[63:0];
  assign n953_o = wishbone_debug_in[64];
  assign n954_o = wishbone_debug_in[65];
  assign n955_o = {n213_o, n212_o, n214_o};
  assign n956_o = {n260_o, n277_o, n261_o};
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n957_q <= n732_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n958_q <= n734_o;
  /* soc.vhdl:490:9  */
  assign n959_o = {n785_o, io_cycle_syscon, n786_o};
  assign n960_o = {n760_o, io_cycle_uart, n761_o};
  assign n961_o = {n844_o, uart0_16550_uart0_wb_ack_o, n842_o};
  /* soc.vhdl:838:13  */
  always @(posedge system_clk)
    n962_q <= uart0_16550_irq_l;
  /* soc.vhdl:838:13  */
  assign n963_o = {n762_o, io_cycle_uart1, n763_o};
  assign n964_o = {1'b0, n848_o, 32'b00000000000000000000000000000000};
  assign n966_o = {n764_o, io_cycle_spi_flash, n767_o, 2'b00, n768_o};
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n967_q <= n714_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n968_q <= n715_o;
  /* soc.vhdl:490:9  */
  assign n969_o = {n775_o, io_cycle_icp, n776_o, n774_o, n773_o};
  assign n970_o = {n781_o, io_cycle_ics, n782_o, n780_o, n779_o};
  assign n971_o = {n901_o, gpio_intr, ext_irq_sdcard, uart1_irq, ext_irq_eth, uart0_irq};
  assign n972_o = {n769_o, io_cycle_gpio, n770_o};
  assign n973_o = {n254_o, n279_o, n255_o};
  /* soc.vhdl:326:9  */
  always @(posedge system_clk)
    n974_q <= n117_o;
  initial
    n974_q = 1'b1;
  /* soc.vhdl:326:9  */
  always @(posedge system_clk)
    n975_q <= rst;
  initial
    n975_q = 1'b1;
  /* soc.vhdl:326:9  */
  always @(posedge system_clk)
    n976_q <= rst;
  initial
    n976_q = 1'b1;
  /* soc.vhdl:326:9  */
  always @(posedge system_clk)
    n977_q <= rst;
  initial
    n977_q = 1'b1;
  /* soc.vhdl:326:9  */
  always @(posedge system_clk)
    n978_q <= rst;
  initial
    n978_q = 1'b1;
  /* soc.vhdl:326:9  */
  always @(posedge system_clk)
    n979_q <= rst;
  initial
    n979_q = 1'b1;
  /* soc.vhdl:326:9  */
  always @(posedge system_clk)
    n980_q <= rst;
  initial
    n980_q = 1'b1;
  /* soc.vhdl:326:9  */
  always @(posedge system_clk)
    n981_q <= rst;
  initial
    n981_q = 1'b1;
  /* soc.vhdl:326:9  */
  always @(posedge system_clk)
    n982_q <= rst;
  initial
    n982_q = 1'b1;
  /* soc.vhdl:326:9  */
  always @(posedge system_clk)
    n983_q <= alt_reset;
  /* soc.vhdl:490:9  */
  assign n984_o = n487_o ? n708_o : current_io_decode;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n985_q <= n984_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n986_q <= n717_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n987_q <= n718_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n988_q <= n719_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n989_q <= n720_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n990_q <= n721_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n991_q <= n722_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n992_q <= n723_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n993_q <= n724_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n994_q <= n725_o;
  /* soc.vhdl:490:9  */
  assign n995_o = {n257_o, n273_o, n258_o};
  assign n996_o = {n783_o, io_cycle_external, n784_o};
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n997_q <= n711_o;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n998_q <= n694_o;
  /* soc.vhdl:490:9  */
  assign n999_o = n492_o ? 1'b0 : n1000_q;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n1000_q <= n999_o;
  /* soc.vhdl:490:9  */
  assign n1001_o = n492_o ? 1'b0 : n1002_q;
  /* soc.vhdl:490:9  */
  always @(posedge system_clk)
    n1002_q <= n1001_o;
endmodule

module microwatt
(
`ifdef USE_POWER_PINS
   inout vccd1,
   inout vssd1,
`endif
   input  ext_clk,
   input  ext_rst,
   input  uart0_rxd,
   input  [3:0] spi_flash_sdat_i,
   input  [31:0] gpio_in,
   input  jtag_tck,
   input  jtag_tdi,
   input  jtag_tms,
   input  jtag_trst,
   input  [7:0] simplebus_bus_in,
   input  simplebus_parity_in,
   input  simplebus_irq,
   input  alt_reset,
   output uart0_txd,
   output spi_flash_cs_n,
   output spi_flash_clk,
   output [3:0] spi_flash_sdat_o,
   output [3:0] spi_flash_sdat_oe,
   output [31:0] gpio_out,
   output [31:0] gpio_dir,
   output jtag_tdo,
   output simplebus_clk,
   output [7:0] simplebus_bus_out,
   output simplebus_parity_out,
   output simplebus_enabled);
  wire system_rst;
  wire [103:0] wb_simplebus_out;
  wire [65:0] wb_simplebus_in;
  wire [28:0] wb_simplebus_adr;
  wire [63:0] wb_simplebus_dat_o;
  wire wb_simplebus_cyc;
  wire wb_simplebus_stb;
  wire [7:0] wb_simplebus_sel;
  wire wb_simplebus_we;
  wire [63:0] wb_simplebus_dat_i;
  wire wb_simplebus_ack;
  wire wb_simplebus_stall;
  wire [68:0] wb_ext_io_in;
  wire [33:0] wb_ext_io_out;
  wire wb_ext_is_simplebus;
  wire [29:0] wb_simplebus_ctrl_adr;
  wire [31:0] wb_simplebus_ctrl_dat_o;
  wire wb_simplebus_ctrl_cyc;
  wire wb_simplebus_ctrl_stb;
  wire [3:0] wb_simplebus_ctrl_sel;
  wire wb_simplebus_ctrl_we;
  wire [31:0] wb_simplebus_ctrl_dat_i;
  wire wb_simplebus_ctrl_ack;
  wire wb_simplebus_ctrl_stall;
  wire n12_o;
  wire n14_o;
  wire [28:0] soc0_wb_dram_in_adr;
  wire [63:0] soc0_wb_dram_in_dat;
  wire [7:0] soc0_wb_dram_in_sel;
  wire soc0_wb_dram_in_cyc;
  wire soc0_wb_dram_in_stb;
  wire soc0_wb_dram_in_we;
  wire [29:0] soc0_wb_ext_io_in_adr;
  wire [31:0] soc0_wb_ext_io_in_dat;
  wire [3:0] soc0_wb_ext_io_in_sel;
  wire soc0_wb_ext_io_in_cyc;
  wire soc0_wb_ext_io_in_stb;
  wire soc0_wb_ext_io_in_we;
  wire soc0_wb_ext_is_dram_csr;
  wire soc0_wb_ext_is_dram_init;
  wire soc0_wb_ext_is_eth;
  wire soc0_wb_ext_is_sdcard;
  wire [31:0] soc0_wishbone_dma_in_dat;
  wire soc0_wishbone_dma_in_ack;
  wire soc0_wishbone_dma_in_stall;
  wire soc0_uart0_txd;
  wire soc0_uart1_txd;
  wire soc0_spi_flash_sck;
  wire soc0_spi_flash_cs_n;
  wire [3:0] soc0_spi_flash_sdat_o;
  wire [3:0] soc0_spi_flash_sdat_oe;
  wire [31:0] soc0_gpio_out;
  wire [31:0] soc0_gpio_dir;
  wire soc0_jtag_tdo;
  wire [103:0] n15_o;
  wire [63:0] n17_o;
  wire n18_o;
  wire n19_o;
  wire [68:0] n20_o;
  wire [31:0] n22_o;
  wire n23_o;
  wire n24_o;
  localparam [68:0] n27_o = 69'b000000000000000000000000000000000000000000000000000000000000000000000;
  wire [29:0] n28_o;
  wire [31:0] n29_o;
  wire [3:0] n30_o;
  wire n31_o;
  wire n32_o;
  wire n33_o;
  localparam n34_o = 1'b0;
  localparam n36_o = 1'b0;
  wire [28:0] n44_o;
  wire [63:0] n45_o;
  wire n46_o;
  wire n47_o;
  wire [7:0] n48_o;
  wire n49_o;
  wire [29:0] n50_o;
  wire [31:0] n51_o;
  wire n52_o;
  wire n53_o;
  wire n54_o;
  wire n55_o;
  wire [3:0] n56_o;
  wire n57_o;
  wire simplebus_0_wb_ack;
  wire simplebus_0_wb_stall;
  wire [63:0] simplebus_0_wb_dat_r;
  wire simplebus_0_wb_ctrl_ack;
  wire simplebus_0_wb_ctrl_stall;
  wire [31:0] simplebus_0_wb_ctrl_dat_r;
  wire simplebus_0_clk_out;
  wire [7:0] simplebus_0_bus_out;
  wire simplebus_0_parity_out;
  wire simplebus_0_enabled;
  wire [65:0] n68_o;
  wire [33:0] n69_o;
  assign uart0_txd = soc0_uart0_txd;
  assign spi_flash_cs_n = soc0_spi_flash_cs_n;
  assign spi_flash_clk = soc0_spi_flash_sck;
  assign spi_flash_sdat_o = soc0_spi_flash_sdat_o;
  assign spi_flash_sdat_oe = soc0_spi_flash_sdat_oe;
  assign gpio_out = soc0_gpio_out;
  assign gpio_dir = soc0_gpio_dir;
  assign jtag_tdo = soc0_jtag_tdo;
  assign simplebus_clk = simplebus_0_clk_out;
  assign simplebus_bus_out = simplebus_0_bus_out;
  assign simplebus_parity_out = simplebus_0_parity_out;
  assign simplebus_enabled = simplebus_0_enabled;
  /* asic/top-asic.vhdl:81:12  */
  assign system_rst = n14_o; // (signal)
  /* asic/top-asic.vhdl:84:12  */
  assign wb_simplebus_out = n15_o; // (signal)
  /* asic/top-asic.vhdl:85:12  */
  assign wb_simplebus_in = n68_o; // (signal)
  /* asic/top-asic.vhdl:88:12  */
  assign wb_simplebus_adr = n44_o; // (signal)
  /* asic/top-asic.vhdl:89:12  */
  assign wb_simplebus_dat_o = n45_o; // (signal)
  /* asic/top-asic.vhdl:90:12  */
  assign wb_simplebus_cyc = n46_o; // (signal)
  /* asic/top-asic.vhdl:91:12  */
  assign wb_simplebus_stb = n47_o; // (signal)
  /* asic/top-asic.vhdl:92:12  */
  assign wb_simplebus_sel = n48_o; // (signal)
  /* asic/top-asic.vhdl:93:12  */
  assign wb_simplebus_we = n49_o; // (signal)
  /* asic/top-asic.vhdl:94:12  */
  assign wb_simplebus_dat_i = simplebus_0_wb_dat_r; // (signal)
  /* asic/top-asic.vhdl:95:12  */
  assign wb_simplebus_ack = simplebus_0_wb_ack; // (signal)
  /* asic/top-asic.vhdl:96:12  */
  assign wb_simplebus_stall = simplebus_0_wb_stall; // (signal)
  /* asic/top-asic.vhdl:99:12  */
  assign wb_ext_io_in = n20_o; // (signal)
  /* asic/top-asic.vhdl:100:12  */
  assign wb_ext_io_out = n69_o; // (signal)
  /* asic/top-asic.vhdl:101:12  */
  assign wb_ext_is_simplebus = soc0_wb_ext_is_dram_csr; // (signal)
  /* asic/top-asic.vhdl:104:12  */
  assign wb_simplebus_ctrl_adr = n50_o; // (signal)
  /* asic/top-asic.vhdl:105:12  */
  assign wb_simplebus_ctrl_dat_o = n51_o; // (signal)
  /* asic/top-asic.vhdl:106:12  */
  assign wb_simplebus_ctrl_cyc = n53_o; // (signal)
  /* asic/top-asic.vhdl:107:12  */
  assign wb_simplebus_ctrl_stb = n55_o; // (signal)
  /* asic/top-asic.vhdl:108:12  */
  assign wb_simplebus_ctrl_sel = n56_o; // (signal)
  /* asic/top-asic.vhdl:109:12  */
  assign wb_simplebus_ctrl_we = n57_o; // (signal)
  /* asic/top-asic.vhdl:110:12  */
  assign wb_simplebus_ctrl_dat_i = simplebus_0_wb_ctrl_dat_r; // (signal)
  /* asic/top-asic.vhdl:111:12  */
  assign wb_simplebus_ctrl_ack = simplebus_0_wb_ctrl_ack; // (signal)
  /* asic/top-asic.vhdl:112:12  */
  assign wb_simplebus_ctrl_stall = simplebus_0_wb_ctrl_stall; // (signal)
  /* asic/top-asic.vhdl:149:19  */
  assign n12_o = ~ext_rst;
  /* asic/top-asic.vhdl:149:31  */
  assign n14_o = 1'b1 ? n12_o : ext_rst;
  /* asic/top-asic.vhdl:152:5  */
  soc_4096_100000000_0_0_4_0_4_0_4_1_4_4_1_2_2_32_529beb193518cdd5546a21170d32ebafc9f9cb89 soc0 (
`ifdef USE_POWER_PINS
    .vccd1(vccd1),
    .vssd1(vssd1),
`endif
    .rst(system_rst),
    .system_clk(ext_clk),
    .wb_dram_out_dat(n17_o),
    .wb_dram_out_ack(n18_o),
    .wb_dram_out_stall(n19_o),
    .wb_ext_io_out_dat(n22_o),
    .wb_ext_io_out_ack(n23_o),
    .wb_ext_io_out_stall(n24_o),
    .wishbone_dma_out_adr(n28_o),
    .wishbone_dma_out_dat(n29_o),
    .wishbone_dma_out_sel(n30_o),
    .wishbone_dma_out_cyc(n31_o),
    .wishbone_dma_out_stb(n32_o),
    .wishbone_dma_out_we(n33_o),
    .ext_irq_eth(simplebus_irq),
    .ext_irq_sdcard(n34_o),
    .uart0_rxd(uart0_rxd),
    .uart1_rxd(n36_o),
    .spi_flash_sdat_i(spi_flash_sdat_i),
    .gpio_in(gpio_in),
    .jtag_tck(jtag_tck),
    .jtag_tdi(jtag_tdi),
    .jtag_tms(jtag_tms),
    .jtag_trst(jtag_trst),
    .alt_reset(alt_reset),
    .wb_dram_in_adr(soc0_wb_dram_in_adr),
    .wb_dram_in_dat(soc0_wb_dram_in_dat),
    .wb_dram_in_sel(soc0_wb_dram_in_sel),
    .wb_dram_in_cyc(soc0_wb_dram_in_cyc),
    .wb_dram_in_stb(soc0_wb_dram_in_stb),
    .wb_dram_in_we(soc0_wb_dram_in_we),
    .wb_ext_io_in_adr(soc0_wb_ext_io_in_adr),
    .wb_ext_io_in_dat(soc0_wb_ext_io_in_dat),
    .wb_ext_io_in_sel(soc0_wb_ext_io_in_sel),
    .wb_ext_io_in_cyc(soc0_wb_ext_io_in_cyc),
    .wb_ext_io_in_stb(soc0_wb_ext_io_in_stb),
    .wb_ext_io_in_we(soc0_wb_ext_io_in_we),
    .wb_ext_is_dram_csr(soc0_wb_ext_is_dram_csr),
    .wb_ext_is_dram_init(),
    .wb_ext_is_eth(),
    .wb_ext_is_sdcard(),
    .wishbone_dma_in_dat(),
    .wishbone_dma_in_ack(),
    .wishbone_dma_in_stall(),
    .uart0_txd(soc0_uart0_txd),
    .uart1_txd(),
    .spi_flash_sck(soc0_spi_flash_sck),
    .spi_flash_cs_n(soc0_spi_flash_cs_n),
    .spi_flash_sdat_o(soc0_spi_flash_sdat_o),
    .spi_flash_sdat_oe(soc0_spi_flash_sdat_oe),
    .gpio_out(soc0_gpio_out),
    .gpio_dir(soc0_gpio_dir),
    .jtag_tdo(soc0_jtag_tdo));
  assign n15_o = {soc0_wb_dram_in_we, soc0_wb_dram_in_stb, soc0_wb_dram_in_cyc, soc0_wb_dram_in_sel, soc0_wb_dram_in_dat, soc0_wb_dram_in_adr};
  assign n17_o = wb_simplebus_in[63:0];
  assign n18_o = wb_simplebus_in[64];
  assign n19_o = wb_simplebus_in[65];
  assign n20_o = {soc0_wb_ext_io_in_we, soc0_wb_ext_io_in_stb, soc0_wb_ext_io_in_cyc, soc0_wb_ext_io_in_sel, soc0_wb_ext_io_in_dat, soc0_wb_ext_io_in_adr};
  assign n22_o = wb_ext_io_out[31:0];
  assign n23_o = wb_ext_io_out[32];
  assign n24_o = wb_ext_io_out[33];
  assign n28_o = n27_o[29:0];
  assign n29_o = n27_o[61:30];
  assign n30_o = n27_o[65:62];
  assign n31_o = n27_o[66];
  assign n32_o = n27_o[67];
  assign n33_o = n27_o[68];
  /* asic/top-asic.vhdl:229:51  */
  assign n44_o = wb_simplebus_out[28:0];
  /* asic/top-asic.vhdl:230:51  */
  assign n45_o = wb_simplebus_out[92:29];
  /* asic/top-asic.vhdl:231:51  */
  assign n46_o = wb_simplebus_out[101];
  /* asic/top-asic.vhdl:232:51  */
  assign n47_o = wb_simplebus_out[102];
  /* asic/top-asic.vhdl:233:51  */
  assign n48_o = wb_simplebus_out[100:93];
  /* asic/top-asic.vhdl:234:51  */
  assign n49_o = wb_simplebus_out[103];
  /* asic/top-asic.vhdl:241:49  */
  assign n50_o = wb_ext_io_in[29:0];
  /* asic/top-asic.vhdl:242:49  */
  assign n51_o = wb_ext_io_in[61:30];
  /* asic/top-asic.vhdl:243:49  */
  assign n52_o = wb_ext_io_in[66];
  /* asic/top-asic.vhdl:243:53  */
  assign n53_o = n52_o & wb_ext_is_simplebus;
  /* asic/top-asic.vhdl:244:49  */
  assign n54_o = wb_ext_io_in[67];
  /* asic/top-asic.vhdl:244:53  */
  assign n55_o = n54_o & wb_ext_is_simplebus;
  /* asic/top-asic.vhdl:245:49  */
  assign n56_o = wb_ext_io_in[65:62];
  /* asic/top-asic.vhdl:246:49  */
  assign n57_o = wb_ext_io_in[68];
  /* asic/top-asic.vhdl:252:9  */
  simplebus_host simplebus_0 (
    .clk(ext_clk),
    .rst(system_rst),
    .wb_cyc(wb_simplebus_cyc),
    .wb_stb(wb_simplebus_stb),
    .wb_we(wb_simplebus_we),
    .wb_adr(wb_simplebus_adr),
    .wb_dat_w(wb_simplebus_dat_o),
    .wb_sel(wb_simplebus_sel),
    .wb_ctrl_cyc(wb_simplebus_ctrl_cyc),
    .wb_ctrl_stb(wb_simplebus_ctrl_stb),
    .wb_ctrl_we(wb_simplebus_ctrl_we),
    .wb_ctrl_adr(wb_simplebus_ctrl_adr),
    .wb_ctrl_dat_w(wb_simplebus_ctrl_dat_o),
    .wb_ctrl_sel(wb_simplebus_ctrl_sel),
    .bus_in(simplebus_bus_in),
    .parity_in(simplebus_parity_in),
    .wb_ack(simplebus_0_wb_ack),
    .wb_stall(simplebus_0_wb_stall),
    .wb_dat_r(simplebus_0_wb_dat_r),
    .wb_ctrl_ack(simplebus_0_wb_ctrl_ack),
    .wb_ctrl_stall(simplebus_0_wb_ctrl_stall),
    .wb_ctrl_dat_r(simplebus_0_wb_ctrl_dat_r),
    .clk_out(simplebus_0_clk_out),
    .bus_out(simplebus_0_bus_out),
    .parity_out(simplebus_0_parity_out),
    .enabled(simplebus_0_enabled));
  assign n68_o = {wb_simplebus_stall, wb_simplebus_ack, wb_simplebus_dat_i};
  assign n69_o = {wb_simplebus_ctrl_stall, wb_simplebus_ctrl_ack, wb_simplebus_ctrl_dat_i};
endmodule

